BSV1       �� BST1   /�zw                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                Compatibility                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                � �                                                                                                                                                                                                                                                                                                                                                                       �                                                                                               " , K . ` � �U                              ��                                                                                                                                                                                                                                                       ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������         S�=|��G                    �           ��� �    �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          ?  08<��_�W+
��I�r�L�c1������m6�]�w�].�[��K%)��U�u��~��g���V�a�x��{��O�S��J���D�a��\�g3��S�T����l+�����h�j����Q�t��v�M&3���i��]��{=�W+�J���`(4���_�W+�J���X&�Y�v���x�w;�N��P�����R	�b������P������I$�y�~���s�\��s9�w���W���U*5-+�J!�h*���f��d)�j
%��t�������m6;�S)�u��~  �x�n�E��x�n�B�@  0�|��w�].7��f	���h��z�N�C�P�d�T
%)*��M��y<�?���q8<>�_/��H��x.7�M&3�����p�l��j��r�L��h�j�J�B�@ ��X�f	�b�r���C��H��x.7���x.7����i��].7�M��y�~�A����������F�A��X�����Z���x��{=���{=��w;�N  0�|�o7�c�X����t-�k��M&3����a����G���T�e����O�S)��U����n�K%�i�������z��s��N���p�l���z���c1,6;'��B�@ �p,�{=���{���g��l+��E"��L��q��^�C���D��H�b�H�b�d�i�z��G��h��z���c1,�{=��k��M&�Y,�{=�o�[-��j�e�y�~���q��^��c���F�����������@�����B�@��P��R�D!���J���`(4���_�W+�e29�n�K�R	�b�H�b�����`(��].7#�d����b��D�P�����R����`�t��v�M���|�o�[��������K����R	"1���K%�i��].�[�V���`����E�q����g�Y�v�F�A�p��V��p,�{�^�G��h������U����n�K������d�i��].�[-+
�R	�b��D���D�P���I$���^�G�Q(�z�g�����e29.7���a0�|��k5��v�����t�m��}>���w;�N�A��X����^  0�|/�K%�i4�}�?�����\'�D���X�s9�n�����T�e2��N���@ ���L����J��p,����_/�K�R�D!��T
���d��t�m6;���c�X���i4�}��_���u���_/��A 0�|�o7��f�I$�y<>?��c1�l�k5��v���S�T
%������S)���j�J����P�d���Z#�d)*5��v��h�u:��O��i4�}>�_����z�g�Y��[�V!�t�V��p��V�B����@ ���L�Q����f����I�r�f	�q�|�W�U��z�S)*5��v��C��H�q8�~��c�X���i��].����[-+�J��A�p�l+��E�q�����s9���k5��v��C���D��p��[-+
�R	�b���B  ��\�g��l�U��z�����^���p��[���e29��{=/�K%��t���[�V�E�q��^��`��T
�R�D���X��y<>�_/���Q(�z��G#���B���H"�������X��y�~�C�P$��|��k�Z�F�����@  ��\��i4�}>�_�W+��E���\'	�q8<>�_����z��s��N  08��_/��e�y<�?����H"�X��S��J�B����@  �x��W+
%)��z��i�z�g3�L���T�e����O�S)�j��E��x��W��j�e29�n�P�d�i4�}����?��g3�L���x.7��f�D!�����b�H��x�n��e29.��m6;�������N  ����G�Q(�z���y<>��o7��C!�h�u:��O'���������A �����c�X����^�@ �p,6;�N��a�����c1������m�{=�W+��E�����G�Q�t��K%�i�����k5-�k5�������m�{�^��c��L��q8<�?�C!�t�V�����T����l�U*��M&3�L#�H��Q�t�m6�]��{�^�G�Q����f�D�a0�|��k5�V���Q(�z����|��w�]��{=��w;'�����P�r�f�D�����F�������@  ���N�A �x�n����P��R	"1��V�E���\��s9.7�c���F�`(�z�S��J���`(4�}>?�O�����M�s�\'����I$29�����z'����I�r��F����D�a�x�n��p,��}�?�G#$29.��m6�������].�[��K�R�D�a08<>��o7����p�l�U*�Z�c1������Y,�{����s9���k5�m����_�����]���}������o7�M�s9.7��f���R	"1,6���W+��r�L����\�g3&3�L��q8�~��a0�|�o�[���e��|/�K��I��Y,6�]���}>?���s�\��s��N���P���l��u�}>?������F��`�h�j�J�a�x.��m6�������].7���S�����Q�t-����]�w;����q�|��w;��s�\�S)�j��E"1��V��b�H��Q(������u:=���u:�^�G��h�j
%�i4��~�O'�I�r�f��B�`�h���j��r���|��k���f��d�i4:=��k��M&3�L�Q�t��v��C!(�z���y�~�A�p��[��������K%)�j�J���X�f�I$��|�W+�e�y<��_/�K%�i��]�w��n�K%�i���n���r���C��H"�X�f����I$29����u�}>?�����|/�K���d��t��v�M&3�L�c�X�f�D�a08<���?�@  0��^�C�P$����O��i�z�N��@ ��X�f�I$2���G#�d��t�V!����f�I�r����a0��^�G�Q�t���[-���z�N�@ �p�v���S��J�B�`(�z��s�\����|/��e2��N�A��X�s9����u:=��w;�g�Y��[��K������d�i��].�[���e29.7����i4�}>?�C!(�z���c1,6����k�Z#�H�q8<>�_/�K�R�D��p���K%)*5��K%�T
%�i4��~�O'�I$��|/��e������s9�n�E���\�����^�A 0�|�o�[-�U*5��K%)�u��~��g3�L�c�X&�Y,�{=/��e29�w�������]��{�^�������G��h�j�J�B��P����d��t�������������m���~�O'�D�a���N ������a�x.7����p,6;��G#�H�b��Y���m6;'�D�a0�����s9�����z��G�Q�t��v��C!�h��U��z��G�Q���M&3���C!��T
%�i�z���y�~�����\'�I����V�B�@����D��H�b��D��H��x�n�P$�y<>?������F���@����D�a0�|/��e2������x�n�E����N�A �x��W�U*�������Z�F  08<��_����z�N��`(4:��O��i4:=/���r&3�f��d��t�m6;����q8<���?���������s9��W+
%����M&�����e29���k5-+����Q��Z��h*��M&3&��l����].7�F��P���l��u����o���v�M�����O'���R	"�����a0��^�C!�h����U*5�m6;��G#�H�b���I$���^�C�P�r�L��q8<>?��g3���C!��T
�R	��Q�t-�U��z���c��L�c��L#�H��Q(�z�N�@  �x�n����Y,����_/�K��I��Y�v�Q��Z��q���O�����M�s��N��`�h�j�J����P����d)�j��E"1��[-+��E"�X���i�z��i��].7�Q�t�m��}>��o7#�r�f	�q8�~����y<��?�O'�I�r��S��J��H�b�r��F�@ ����F�@���H�b�d�i4:������|��w�]�w;�N�A�p��V�B��@��P�d)�j����Q(4����o7�F��@  08����w�].7�M�s9�w��n��e29����u:�����y�~��g3�L�c�X�f����`�h*5��v��q�|��w�].7�c1����e2���G����J!(4:��O��i4:�^���P��Y�������v��f��B��@ ���L�Q(4�}>���w;���������y�~����y�~��c�X�f�I$���^���q��^�G#�r�L��q8<>�_/��e29��{�������^�����D�����F�`�h�j�J��A ����G#���I$��|�o7�Q(4:�^�G�Q(4:��O����Z�F���P$��|��w;�N�`(�z�N�C��H"�X&��l+
%�i�z�N�C!(4��~��a08�~�O�S�T�����V�B �p,�����o�[�V�B  �x�n�B�@�`��Z��h�j�e��|���{�^��a0��^�C��H��Q(�z'�I$�y���o7�M�s���G�Q(�z���c��L��q8�~�O'	�b�H�b$2�\��s����c1�l�����U*�Z�F����H��Q(�z��G#�r���C!���J�B��@������A�p�l+����l�U*5�V�E"��L#����V��b�H"���F��`�h*5�V�E�q8<��_/��H��Q�t�V�E��x�n�K%���E�q8<��������_����z'�����d��t-��������u:�^��c����C!�h*5�m6�].��m6;�N��`���J��A�p,6����k�Z�c1,���~���q8�~�O���t��K%�i4���_/��e29�w�].7�Q��Z���a08����w�].7��f	"�X��y�~�O'�����d�T�e2�\��s9�w;�g�����e��|/�a�x.�[���e�y�~�O'��d��J!�h�j
%��J�P�d)�j
�R�D!����E�����G�Q(��].7����\�g�Y������m��}>?�����|��w;�N�C�P�d�i4���_/�K�R	"����C��H"�X&3�L��q8<���?���s9.7�F���H"��L�c�X&�Y�v�M��y�~�G#�H��Q��Z��C!�h�j����l��u:��O�S)��U*5�����v��f�D��p�v������L����J�B�@  0�|�W�U����n���Q(���n����L�c��L#��D��H���h��U��z�g�Y�v���S)*5�m�{�^�������C�P$��|/�K%���Z��q8���o7��C�P�d�T�e29.��m�{=�W����j
�R�D���D���X�f��d)���j��E"1�l��u��~�O'	�q�|/�K%���Z#��R�D��p������m6��n�E"1������m�{�^  0�|��k�Z�c�X�f	�����G�Q(�z��i4:����s�\��s9����u:�^�C!��T
%��J!�h*5��v������Z�c1��[�V�E����N�C!��Z�c1��V�B��P��R�D�����A�p�v�M���|��w;�g�Y,6��n�E�q���O���t����m6�].7�M���|/�E�q8<�?��c1��V�E"�����a08<>�_��k��M&3�f�I$2���G#�H�q���O�S�T
�R�����P�d��t-����]���}�?���q8���o���v#�d)�u�}���������������_/�����T
%��J��A�p,�{�^�G#�H"���F�`��Z���x.7�M�s�\��s9�n�K%����b��D�a�����c1�l�k5�V����h�j��E�q�|�W����j
���d�T
%������S)�j�e�y�~����H�q8�~����y<>�������_/��e2�\�S)�j
�R	�b�d)�j���b���l+���b$2�\'���A 08<>?�O'��B�@ ���L���x.7��C!��T��r&3�L�Q��Z�c1����e�����g�Y�v���a��\��s�\������O�S�T�e�����g��l�U��z�N�C�P$���^��a0�|/���r������X�f��d)�u:���g�Y,���~���s����c1�l�U*�����i�z'	�b�r&3�������L��q�����s���G���T
%�T
����R	��Q(4���_/���r&��l+��E���\������f����I$29�n���Q��Z�c1�v#�H���\���t-�k5��v�F�`�h��U*�Z�F���P�r���C!�h��z�g��l+��E�q8�~�O���t-+�����h�������j������T�e�y��_��k������t�m����������_�W����j��E�q��^�G#�r�f�I�r��F����@ ��X�f�I$29��W�U*5-�k5��v��f��B���@�`��T�e2���G#��D��p����v�c1��[��K%�i�z�S)��U���]�w;��G�Q(4:=�W+�J���D�P��R�D��������p���m6;�g�Y,�{�^��c1�l����j�J�B�@��P��R	��Q(4:=����}����?���q8��_/������V��H����T
%�i�z�N�C!���M&3�f�������I�r���|�W���U����n�E"1,����_��k��M&3�f���A 0�|�W+�e29��W�U��z�N��a0�|�o��m�{=��������k5�m��}>�_/��e2�\�S)*5���e29.�[-��u���_/���X&3�L#�d�i�z�N�C��H"��L���x����u�}��_/����h�u:�^�C!(4�}��_/�������E"1��[���e29����u�}��������o7�M&3�L��q8<���o��m6;����Z�F��`��T
%�i�z�g�Y,6;��s�\'�I$��|��w���W�U�u�}������_��k5�m�{=/��e��|��w;�S��J���`�t�V���`�h���].7���S�T
%��t�m6�]�w�]�w;��G���T
%�T
%��t�m�{=/����h*�Z�F��`���J����B ���L#�H���h*5���e2�\�g3��S)�j���b�r&��l�U*���f�D!�h�j�e����O'�I$2�\��s9��W��j���Y�v��C��H��Q����f�������D���X�����Z�F��@�`��T�e�y<>�_/����P�d)���j���b�H��Q��Z�F��P�d�T��r�s9.7�M&3��F��`��T
%��������J�B  ���N�A 0��^�G#���B��@  08�~���s��N�������C��H�b��D!��T��r����a�x�n�E"1�l����].7�M�s9��W�����U*5��v��������f	��Q�t�V�����F���P��R��B  ��\'��d)�j���Y��[-�U��z�N�A 08��_/��b�d��J���D��p�v#$���^�A�p,6��n��e�y<>���w�]����~�����|�o�[�V�a�x�n���r�L�c1,�{���g3��S��J�a���N���������p,�{=�o7���x.7�F  0�|/��e2�\�S���E���\��i�z����|���{�^��a�x.7��f�D!�t��v���S)�u�}��?�G�Q(���n���Q��Z�F�A�����C�P�r���|/�E"1,�{=�W+�J���`(4������{�����y�����{�����y��_�W��j��E"1�l���U�u�}�����o7�c1,6��n�E"1�v��q8��_/���r��S)����U����n�E�q��^�G�Q(4��~�O������f�D��p�l��j��E�q�|�W+
����R��B�@  �x��W+�J������������D�a���N���P�d��t�����v��C!��T
����������R�����P���I�����K�R	��Q��Z#$2�\'���R	���h���].7�F���P$��|�W�U*�������Z��C�P�d�i4:�^�����@�`�h��z��G#�r�f���R�D�a08<�?�`(�z��G����J�P�r�s9���k�Z�c�X�����Z�F��@  08<����?�O�S)����n��e2�\�g3�L#�d)��U�u����o7#$29.�[�������V�a�x���k5-+���Y,6;�N��@�`���J���`(4:��O��i��].�[�V�a���N�C!�h�u:=��w�]��{�^��`�t��v�Q(�z���y�~�C�P$29�n�K%��J���`����E"���F������@  0��^�G#$29.�[-��j�������e2��N�@ ��X�f�I$29.7�F�@������A����F�@��P�r�L�Q�t���[��K%�i��].7��f�I������e2��N �p���K%�����Q(�z��G��h�j�e����O���t�m6���W+�J��A�p�l��u:�^�G#�r&3��F����D����L�c��L����\'��d)��U*�Z#��R�D�a�x�n��������e�y�~���s9�n�P�d�T
�R�����P��R����`(4�}��?�O�S�T
��I�r��S)�u:=/�E�q�|��������k���f�I$�y<�����_/�K��I��Y,6;�S)��U*5�m6;�N���P���I�r���i4:=����}�?��g�Y�����[-�����U�u:=/�K���d��t���[����r�L#$2�\�g3��S)���j�J!�t���[�V�B�@�`��T
%�T
%)�����j
��I�r�L��q��^����x���}>?���s9�n����P$��|��k��M���������|�W�U*5�V��b��D!�h��U�u:=/�P��R��B���H�b�r�L�c�X&����K��I$�y��_�W+�J����P$�y��_��k5���e29����u��~�G#�H��x��W+
%����M�s9���k��M�s9.�[��K����������R	"��L��q8���o��m6��n�K%�i4:�^�C!����E"�X��S)�u:=�o��m�{�^��������c�X�s���G#��D!��Z�F  �x��W�U���]����~�G���T�e�y��_/�E"1�l�k���f���A 0�|�o�[-+��E"1,��}>?�O'���A 0���O�S)�j�J����P�r�L���T
%��t-+
��I$�y<��?�G�Q�t-���z��s9.7�Q�t����m���~�O'��B �p������Y,6;'��B��@�`(4:����s9���k5�����Y�v��q�|�o���v���x���}>?�O'�����d��t��v�M���|�W+�e���^�G�����E"1�v�F�A�p,�{=��w;'�I$29.7�M��y<>�_/�E�q8<>�_/��e2�\'�D��H�b���l+
%�i����W��j���Y��[�V!(�z�g��l��j�J�a�x�n�K%����M&��l�k5��v�F�A�������p��[-��j
%)��U*���f	��x�n�B�`��T��������r�L#�H��Q���M����^�A�p�v�F�@�`��T
�R���A��X�s�\�g3���C�P��Y��[���e�y�~�O�����M&3�f�I$2��N���P����V�B �p,�{�^�A �x��W�U*�Z#$�����g3&3����t�V���X�s9�w��n��A �x�n�E�q8<����?��`�t��v�M�s9�n������`��Z�F�����D!�h�u:=/���Q���M&3��F��`����E�q��^���q�|��w�].��m�{=�o���v�M&��l�k5����m�{=�W+�J�a��\�g��l+�J��p,6;'���A ���N�C�P$�y����w;�������N������F���P�r��S��J��A��X�f�I��Y,6�].�[-�U�u:=�o7�c�X�f	����N����H����T�e29�w;�N�A�p��V�a08<����_��k������t��v������Z��q8�~���@ ����F�A �x.7��h��������U����n�K%���Z#��Y,6;���c1��V�E"��L���x�n�K��I$�y<��_�W+���b�r�s9����u�}���_/�a��\�g3�f��d)��U*�Z#���B��@ �p�l��u:=���{=�o��m��}��?��a�x��W+��r&����K%��t���[�V�E�q��^�G#���B  �x�n���Q(��]����~���s��N����X��y<��_/�K%�i��]��{�^��@�`(4:�^��c��L�c����C������`��Z��C!����f��d�T
�R�D�a�x�n��������e29���k5-�U���]��{=/�K%�i�z'����I�r�L�c���F  �x.7���S�T�e�y<�����o7����p�l�k5�m�{���g3������X���i4�}������?��g�����e2���G�Q���M���|��w�]�w;�N�C!(4:=����}�?��`�h��z���������y<>��o��m��}������_���u:��O��i4:=��w��n�P�r�L#�d��J�B�@ ��X���i��]������o7�M&3��S)�j�J���`��Z���a08<>��o7�M&3�L���x�n�K��I�r��F�@ ��X��������y�~�����|����}����w��n�E"��L���T
������d�����f��d�i4:=/�K%�i�����k5-���z�N�A 08<>���w;'������R	�b��Y��[-��u��~�O��i�z�N�A ���N��`(��]��{��O'�������D�����F��`�h�j��E��x��W+���b��D!�h���].�[�V�E��x.7#$2�\�g���V��H���h�j�J��p��V!�h�j�J�a�x.�[�V���D���������X�f��B�@�`(4:=�o7�Q(�z�N��a���N�C!���M&3�L��q8�~�O'	"����C!(4��~����y�~������F�`�h*�Z�F����@ ���L#$��|�o7���S)*5�����v����������������\��s9.7���S���E"��L�Q��Z�c1,����_/������J�a0�|�o7�c1�v�F���P��Y�v��f	"1�v#�H���h�j
%����b��D��H�b$29.7��h�u:=/�K%)�u:�^�G#�H���h�j�J��A �����c1�l��u:�^��`�h��U*��M&��l����]�w�]�w�]����~��g�Y�v��f���R	�b���I$���^��@�`(�z���c�X��y��_/�E"�X��S���E�q��^�@ ��X���i��].�[-+�e�y<>��o�[��K�R�D!�������t�m�{�����y������}���o��m�{�^�`�t�V��b�H�b�H�q8��_/���Q��Z����\���y<>?�C�P��Y��[-��u�}�?��`�h��U�u�}�?��g3��y�~�O'��B ���L��q8�~���s��N�C!�h�j�e29�n��e�y���o7���S)�j
�R	"�����a08���o7����i4���_/��H�b��D�P�r��F�A�p�v���S)�j���b�H�����G���T
%�i4�}��?�O��i4��~���q8�~����x����~�G#��Y,6�].7����p,���~���s9.�[���e29���k5�m6��n�K��I$29���k5-+��r�L�c1��V�B��@  ��\�g�Y,6;����q8<�?�O�S��J���X�s9�w���W�U*��M��y��_��k��M&��l+�����V���X�f	��Q���M��y<��_/�E�q8<������o7#$2�\���t-����]��{��O'��d���Z�F���P�d)��U*5��K%�����Q(�z�N�C�P���l�U��z�g3�����p��V���Q����f	�q�|�o�[���e2��N�����L#�d��t���[�V�a08��_���u:=����z��s�\�g�Y,6;�g3�f�I$�y<��������w�].7#�d�i4�}�?����x.7�c1���m�{=�����]�w�]�w��n�K%�T
�R��B��P���l����j����Q����f���A �x��W+��r�L����\'��B  0�|�����~�O�S����b�����R��B  08��_��k�Z#�H�b���B��@ ����F��`�h�j
%)��z�����x�w;�����x�n��p�l�k5�V�P�d�T
%)����n�K%������S�T
%���E�q8��_�W+�e29����u�����w��n��b��R��B�@��P��R	��Q�t��K�R	�b��Y,6;�N���p�v�M&3&�Y,6�]��{=�o7�M���|/�K%�i4:�^�@ �p�v�F  0�|/�E"�X&3�f���R��B ��X&�Y,6;�S)������k5-+���b�d)�j�e�y�~���P����d��t�����Y�v��f��d�i�z'���R	��x�n���r�L�����N�C!�h����n�B�@  ��\'�I�r�������f����I$�y<>?�O'��d)�j
%��t��v�c1�l�k�Z��C!������Q(4:=����}�?�O'�I$29.7�F�@�`���M&3��F��`�����b��D�P��Y,6�].������v��f�I$�y�~��a�x.��m�{��O�S)*5����m�{�^��c1,6������z�����^���p��[���e2����c1,��}>�_�W+
��I$�y�~���s9��W���U�u:��O�S�T����l�k��������M�s��N ����F�@�`(�z'	��Q(4��~�O'	���\����Z#��D��H"��L��q8<���_/����Y,6������z'�I�������r&3����a08<>?�O���t�������m�{=�o7��f��d��t-�U������k5�m6;�N���@  �x��W�U�u�}>?����y�~�G#���B �p��V�E"�X�s���G�Q��Z���a0��^�G#�����`�t��v�c1��V����L��q8<������{�^�����\�S��J���X�f�I�r�L#��D�a0�|��w�]��{=��w;�N�A �x��W��j�J�B��P$�y���o�[��K�R�D���X�s�\�g��l�����n�K�R�D��H�b�r�L�c1�l��u���_�W+��r�L�c1,6;�N��`�h��U*�����i�����k���f�D!���M��y<>?�G��������h�u��~�G�Q(����W����j��r�L�������c����C��H"1�l����].7�����t������[�V��b�H�q8��_�W+�e�y<���?�O'�I�����K%�T
����R	�b����d�i4����o7��f���R	�q���O���t�m6;����Z���a08���o�[-�k5�V�B��@  �x.���v��f�I$29.��m��}�?��g3�f�I$�y<�?�O'��B��@ ��X�f�D�a�x����u:=��w;�N��a08<>? �p��V�E"1,6�]�w;����q8�~���s9�n�K��I��Y�v#�H��Q(�z��G�Q(��].7���a�x��W������j��E��x��W��j�J��p,6�]���}���_�������W�U*5�m6;�N����H����T����l��j�J��A��X���i�z���c�X�f�I$��|/�E"1���K�R�D���X&3��S�T
%)��U*��M���|/!��T
%��t��v�M&�Y,6��n�a08�~�@�������`�h���]���}>��o7�F���P$2�\����|/�E���\��s9����u�}>?��g3��S)�u:=�������W�U�u:�^�G�Q(4��~�O��i�z�S)�u:=�o7���S)*5-�k���f�I��Y�v���a�x�n�a��\���y<>?�G���T
%��J��p,���~��g3��S)���j�J�B�@  ��\'�D�a0�����s��N�C�������P�d���Z�F��`��Z#��D!�h�j�J��H���\�g3�L#��R������H"�X&3��F�@����D�P�d���E�q�|�o7��q8��_/����Y���m6��n�K�R	���\���y��_/���r��S�T
�R�D�P������I��Y,6;��s9.�����m6;�N��a08<>�_���u:�^�G���T�e����O�S��J�a�x�w�].7�M���|/��A�p��V��A�p,6;�N��P$��|������_��k5�m6;��i����W�U����n�K%�i�z��G#�d)��z�N�A �x.�[-��u������{����s9�n�K���d�T
%��t�V�E������c1��V���`����������E�q8<�����?�O'�I$2��N�C��H�����G#��R�D��p�l���z�g3&�Y���m�{��O�����M��y����w����k5�m6;�S)�j���b�d)*5-�k�Z#��D��H���h*�Z�c1��[-���z�g3����a��\�S�T
�R	��Q(�z����Z���a����G�Q(��]���}���?�O'��d���E�q8<>?�O�S)������k5-�k��M&���V�B�@  �x���k5��K��I$�y<>?�O����Z�Q���M&3�L�c�X&3�f����I�r�f	�b�H�����J�B  �x����~��c��L�Q�t�m6���W����j
%)*�Z���a�x�n��e���^��������c���F�A ��������\��������s9���}>���w;�N��a08<>���w;�N�A ��\�g3�L�c�����a���N�C��H�b�r�L��h*�Z�����X�f	����T���Y����v��C!�t���[-��u:�^�A 0��^�G��h����n���X&3�������f���A ���N��a08��_�W+
%�i4:=�o7#���l��u:=��k5��K%���Z�c1��[-�k5�����Y,��}��������w;�N���p,6�].�[-+�����V�B�@��P$29��W��j�J�B��P$�y��_�W�U�u�}>?�����|��w;��G#�d����M&3&3��S)�j��E"1���K�R�D���X&3�f����I$2�\�S��J�a08�~���s��N���@  0��^�G#�H�b�r&3�L��������h�j�e��|�W+
���d�i��]��{�^���p���K%�T
%)�����j��E"1�����r�f�����P�d�i4:�^�@  ��\'�I$2�\�g3���C�P�d��t�m6;'	�b�d������S����b��D�P��R��B����@�����B �p,6����������k�Z#$29.�[-��u�}���������_/�����l�U����n������C!�����b���I$�y<>?�G�Q��Z�Q(�z�g�Y����v�c1���K%���Z�Q��Z�c1�v�F �p������Y����v#��D��p�l��u�}���_�W�U�u:��O��i4�}>?���P�r�f��B�@ �p���K%)�u�}��_�W�U�u�}>�_�W+
�R����`�h�u:=�W+�e2�\��s��N��a0��^��a08<>?�O'�������D!�h��z��G#�r��F ����F�@����D�a0�|��w�]�w�]�w;�N���p,��}>������~�O'��d�i����W�U*5�V����h�u��~�G��h���j�����h�u�}>���w;'�D�a0�|/�B��@ �p��V��H�b$29.�[�V���X�f����I$29.�[-�k����S)�j�J�B��@�`�h*��M&�Y,�{�^���p�l�k�Z�F������@�`(4:=/�B�@�`����f	�b�d�i���n��e�y<�?��g3�s�\��s9�n���Q(4:=/�K�R	���\���y��_�����]�w;�g��l��u�}���_/��e���^��c1�v����i4:=/�E"��L��h*5���[����r�s9.��m�{=���u��~��P�d�T
��I�r��F��P�d�i�z�����^����X��y<>�_/��e2�\�g����K�R�D!��T��r�L��q����g�Y���m�{=�o�[-+�J���X���|�o7�����t�m�{��O'�I�r��y�~�C!�t������[��K�R����`�t-�k5�m����_��k5���[-+��E��x�n��A 0�|/������V�B �p,������w;�N��a0�|/��e���^���q8�~�G�����E"1����v���S)�u��~�G#�d)*�Z#�H��Q(4��~�A�p��[-�k�Z��C!(���n����Y,6;���c1�v���S)����U*�Z�c�X����^��a��\����|�o�[�V��p�l��u�}>?�A������a�x�w;�N��`�t��K%��t��v���a���N�C��H��x��{=/��A 08<>�_/������������J���`�h��U*���f	"1��V�E�q��^�G��h*5�m6��n�K%��t-�������k5�V�����T
�R����`�t-��j��E"�X�f�I$�y<��������~�O�S�T��r��F��@  �x.�[-���z�S)�j�J����L��q�|������_�W�U*5���[-��u�}��?�C�P�d)*5�V��p��V��b�H�b�r�f	����N�C!�h*5��v�M�s9.7�F�A ���N���p��V�B�@�`�t���e2�\����Z�c�����a�x���k5�m6��n�E�q��^����x���k����S�T
%�i4:=�o7�F�A�p�l+�J!�h�u���_�W���U*5��v����i4:�^�G�Q�t�m��}������?�O��i4:�^�G��h��z���y<>��o7���S)���j��E"1,����_/�B�@�`��Z�F�`�h�u:���g�����e�y<�?��a0�|�o7�F  08�����{�^�G#��D�a08<>���w;�N��a�x����u:=�o7�M&�Y�v�F  08�~������B��P$2�\����Z��C�P�r�L���x�w;'��B�`�h��U*5�m������������w��n�������E���\�����^���P�d���Z��C!(4���_���u:=��w�]��{��O�S)*�Z����p�l�U�u�}���_�W�U�u���_/�P$�y��_/�E"��L#�H��Q�t�m�{=��w�]��{=��k�Z�Q(4��~�O�S��J�B��@����D��p,�{���g����K%����M&��l+�J�B���@�`���M��y<>�_��k��M&3�L���T��r��F�A���L#����d�i��]�w;����|/�K%�i��].7���x�����z'���R���A 0�|�o7�M�s��N �������p�l+����Q(4:=�W+��E��x�n�K��I$�y<>?���s9��W���U*�Z�F�`���J������C!����E"1�v������G#�H��Q(�z�N�C!�����b���B  08<��_������n���Q(4:��O���t-��u�}>������~�A�p���K%�T
%��t����m�{=�o7�M&3���C�����A�p��V��b�d���Z��C�P�r�L��q�|���{=/�K%��t-�k�Z�c�X��y�~���q���O'���R	�b��R	���h�j�J��p����v�F����H����N��a0�|����z�N�C!�h��z'�I$��|�o�[��K�R	�q8���o7��h����U*5�m����_/�E�q��^�G#�����������`�h*�Z�F�A �x��W��j�e29�w;��s9.7����i4:�����y<>���w;'�I���l��u�}��_�W+
�R���A ��\'	�q8�~����X�f	"�X��S����b�H�b�d���Z������L�Q(�z���y<>?��g����K%)���j
�R	����T���Y��[-���z�g3�f�D��p��V�E�q��^�A��X&���V!(����W��j�J��A���L#�d�i4:����s�\'�I�r�f����`��T
%�i4:�^�@  08<���?����x.7�Q�t�V�E�q8���o7#�H��Q�t�V�E"1�l��j���b��D!�����b$�y<����w;��i4:��O�������S)*5���e2��������N����X&�Y�v��q8<>?�O��i4:=�o7���S�T
�R�D��H"1�����[��K��I�r��F  08����w;���c�X�s9.7��C!(4����o�[-�k5��v��f����`(�z��i4:�^��c1����e����O'���R	"1,�{�^���q�|��w;�S���E"1�l����j�J!�h���j�J��H�b��R	�b����d�i4:��O'����I������e29.7��C!��Z�F�A 08<>?����x�w��n�B�@ ���L�c���F�A����F�`�t-�������k5�m6���W+���b����d����������M&�Y,�{=�W+
%�T����l��u:�^�C�����A ��\��s��N�C!��T
�R�������D�a�x.7���S�T
%)*5�m�{�^�G#$29��W���U����������n���r��S��J�B�`�h�j�J�B���@ ��X�s9����u���������_�W+��E"1�l��u����o7�F�A �����c��L#�r��y��_���u���_��k�����i���n!(���n��e2�����q8�~��g�Y����v�M��y<>���w;��G#��D�a0��^���p�l+�e�y�~���s9�n�K%�i��]��{=�o���v�������M&3&3�f�I$�y<>�_���u�����w�]����~�����|������_/�a�x.���v�M�s�\'�D��H���h��z�N����@�`���J�B��@��P��R	�q��^�A 08<�?�O'�I$2�����q8�������~�O'�D��p��V�����H"1,6�].7���S���E"���F �����C!�h��z�N�A�p,�{=�o7�c1�v��f��d)�j��E"1,6�]�w�]�����_/���r��S���E�������q8<>?���s�\'�D�a�x�n��e�y�~�O�S)�j
%������S��J��A�����C�P��R�D�a��\��s9��������{=���u�}�?������B�@���H"1��V�B���H"��L�c��L�c1,6;'�����d�i4�}>��o7���S���E"�X��y<>��o����[-�k5-+
�R	"1�l�k5���[��K��I$������s�������\'�I���l+�J��A ��\���y�~��c1��������[��K��I$29�w;�����^�C�P$��|�o�[�V�E"����C�����A�p�����r�L#��D���D�a08�~���q�|�o��m������w;�����M������g��l��u��~����H���\��i���n����L���x�n��b���B�`(��]��{��O'��d������S��J�B�`��T�e29���k�Z������L�c���F�A����F�@ �p,��}�?�O�S)*�Z���x�����z�N�C!�h���j�e�y<��_��k��M&3�L�c1,6;���c1�l+�J�B�`�h�j��E"1�l�k5���e�y�~�C!���J�B  0�|�W+
�R���A�p,������w�].7�M&3��S)�u����o������v��f	��Q(���n��e�y��_/�E"1���K�R�D!(�z�N�������C!�t-���z����q��^��c�X�f��d��J����B����@ �p�l��j�e2���G�Q��Z�c��L���x����~�O'�����d)*�Z�F�A �x.7��f�I�r&�Y,6��n��e29���}����o7�F���H��Q(4:=�o7�M&3��S)��U�u:=������_�W��j��E�q�|�o�[������l���z�����^���q�|/�B����D!(4��~�C�P$29.7���S�����Q(�z'�D���X�s9�n��e�y<>��o7��C����B���@�`�h�u:�^�G�Q(4:����s�\'�I$29�w�].��m6;��G#$2��N��P��R�D�P$29.��m6;�g3������X����^�G��h*5���e��|�W�U*5�m6���W+��r�s9��W+��E"��L�c1����e29.7�M&3���i4�}>������~��g3�L�c�����a���N����@ �p��V�E"1�l+��E"1��V���X��S)���j���b���B  �x.7�F�@�`(4��~��g3�L�Q(���n��b$2��N���@��P�����K�R�D�a08�~�C��H�q��^��c1�v���S)�j
%��t-�k5-+
%��J�B  ��\�g3�s�\�S��J�B���H�q��^�C!��Z�c��L#��D!���M&���V�a08�~��c�X�f�D��p��[-�U�u�}����w�].7��f�I$��������|�W+��r&3���i���n�K��I��Y,����_�W���U��z��G�Q�t�m6����k�Z#�H���\'�I���l+�e29��{=�o7�c1�v�M&�Y�v���x�n����Y,�{�^��c�X�s9���}�������~��`��T
%�i4:����s��N��a0����g3�������s��N�`�t��K�R	����N�A�p����v�M����^�`���J!(��]���}>�_�W�U��z�g3�L�c1�l+
%���Z�c���F���P��R	"�X&3��F�@�`(�z�N�A ���������N�C�P�d��t���[-+�J�B��@�`������i���n����h�j���Y���m6������z�N���p,6;���c�X�f���R	��x�n���r�L��q��^�C�P�d��t-��j�J!�h�������j
�R	�b��R	��Q�t��v��f�I����V��A ����G�Q(����������W�U*����S�T
%)*�Z�c1�l+�J���`��Z��q8�~��g�Y��[-�U�u:=��w;��i�z�N��a��\�S)��U*�Z����p�l��u��~�O�S)*�Z�����X&3&3��F�A��X&�Y�v�M&3��S��J�P$�y<>?����y<��?��c��L�c���F�A��X�s9��W+�e������s�\�g3�L�c1�l�U*�Z��q8��_/�E"1,�{=�o7�����N�����L�c1,�{=/��A ���N�C!�t�m�{=/�P��Y,6;��G#�����`(��].����[�V�E���\�g3�L#�H��x��{�^���p����e��|�o�[-��u���_/���r�L�����N�C�P�d�i4:=���������{=���{=�W����j�����h�u���_��k�Z��C!��T
�R	�b$2��N���P$���^��c1,���~�G#��D��p����v��q�|��k5�m��}>?��@ ��X�f	"��L���T
%)�u��~��������g3��y���o7�����X��S���E�q�����s9��W�������U�u:=/��p����v�M��y<>?�G#$29��W+�J�B�@ �p�l+����Q(�z�N���H���\'�����P�d�T
�R���A ���N��a��\'��d������S)�j�J�a0�����s9�n�K%)��U�u����o7�F��`(4:����s�\�g��l�k5�����v�M&3�L�c�X������g3�L���T
��I����V��A 08�~�G�Q�t�m��}��?�@  0�|/��b�H�b$29�n���r������X�f�I$�y<������}>?�C���D�a0�|�����~�G��h�u:=�o7�M�s����c��L��q���O����Z�F���P$�y���o7����i4:=/�E"1��V��b����A 0�|/�E�q�|�o7��f���A �x�n�B�@�`��T
���d�i�z����|�o�[�V���Q(4:�^��c1�v�M�s�\�S��J�B����D�P�d�i�������z�N���P��R	�q8<��_/�K%��t��K�R	�b�r�f�D!��T
%������S)���]���}>?�G��h��U������k5-��u:=�o���v�F  08����w;�S�����Q�t-+�����V�����F�A��X&�Y,6;���c���F�A�p�l�k5�m�{���g��l�k��M�����O�S�T�e�y<�?����x��{=�o�[�V�a�x��W��j
%�i�z�N��`��T
%�T
%)*�Z�F��`(��].�[-+�J���`�t��K%������S����b�H"1���m��}>?��g��l+����l�U*5����m6;���c�����a0�|/����Y,6;'����I$����O���t-���z��i��]�w;'�I$��|�o7���S�T
%�T
%���Z�F����H"1����e2���G#��D�a��\��s�\����|������_�W��j����l���z�N�C�P$�y�~��g3�L#�H�b���l��u:�^�G�Q(4���_/�B�@�`�h������k5��v��f�I���l����]���}>?�G��h��z��G�Q(��].�[�V��b�H�b���B�`��T
��I�r�L�Q���M�s9�w;'��d��J�B��P$�y�~��g�Y�v��q��^�C!����E��x�w;�N��`(4��~��c1,6�]�w;�g3��S)�����j
��I$����O�����M�s������������x��W+�e29�n���Q(�z�g3�L�����E��x�w��n��e���^���q�|/���X&3�����p��V���`���M��y�~���q��^������F����H��x�w;��G�Q(4:�^��c1�v#$29�w;��G#�H�q��^����@ ��X&3�L�Q(�z����q����g�Y�v�M&3������X�s9.�[���e29��W+��E"���F  0�|��w;��s9�n�����T�e2�\�S)�u��~�������G��h�u�}>�_/���Q��Z��C!��T��r��F �p����e29.�[-+
�R	��Q(�z�N�`(�z��G��h�j
%�i�z�S�T
�R�D�a�x.�[����r�����Z��q��^�G��h��z���y�~�O'�I�r��S)�j�e��|�W�U���].7���S�T����l��u�}>�_/�K%���Z�����X�s�����q��^�A ����G#���B��P���I$��|/�E"1,��}>���w;'���R	"�X��S��J�B�`�h�u�}�?�@  ���N�@���H"����C�P$2��N�A�p�l��u:�^�@�`���J�a0�|�o7��q8<>��o7�M&�Y,6���W���U*5-�U�u:�����y<>?�G�Q�t�m����_/�E"��L#�H"1���K%�i4:=�W�U�u:���g3��S���E"1�v#�r�L#�H�����J�B����@ ����F�A �x�w�].7�Q(4�}>��o7��f	"1�l+��r��S)���j�J�B�`������i4�}>�_���u��~�O�S)�j���b��D���X�f	"1���K%�T
%�����f	"1����e�y<�?�G�Q(4����o7����i�z�S�T��r��F�`�h��z���t�m�����o�[-�k5�V���Q(4:��O��i�z�N����X&��l�k�Z�Q(4��~�O'���R���A�p��[���e29�n���r���|/���X��S)*��M&3��F��@�`��T�e���^�G���T���Y�����[�V��b�H"�����a0����g3�L��q�|�W��j
���d������h���j�J��p���m6���W��j
%���Z����p�l+��E"�X���|�o7���S�T
%�i��].�[-�U�u:=/����h*��M&3��F�@���H"���F�A�p�l+�J�a��\'��d��t-�k5�V�B���H"��L#�r��S)�j
�R	�b�H�b$�y�~��@���H�b�H"���F��P�r��y�~�O'��d)�j
%�T
���d�T
�R�D�a0��^��a08<>���w��n���r���������C��H�q�|/�K�R��B  0�|�o7���S�T
%�i�z�N��P�d���Z��q�|�W+�J�B ����F�A�p,6;��G�Q�t��v�M�s��N�A ��\�������g3�����O'	�q8�~��c1�l�k5�m6;'	�b�d)��U���]�w��n�K��I��Y�v��q8���o7��h�����W+���b��D!(�z��s���G#���l�U�u��~��g����K%���E�q�|�o7�c���F�A����F�`�h���j�J�B��@ �p���m�{��O'����I$29�n�K%�i�z��s�\�S)��z�N�C!�����b�H��x.7�c1�v�c��L#���l��u��~�G#����d��������t�m6�]�w;�S)*5��v���x�����_/!��T�e2�\�S)�j��r�f���A 08�~�G#�H"��L��q��^�G#�d���E"1�l�k�Z#�H�q8<>�_/�K�R	"1���m���~�O��i4:�^�G#�H"����C���D�P�d����M�s�\'��d�i�z'��B�`����E"�X�s9�w;�S�T��r�s9�w����k���f	"�����a�x.��m�{=����}>?���q8<������������o7��f�D��H�b���I��Y�v�F��`��T
�R������H�b�H�b$29��W+��E�q�|�W+�J������C��H��Q(4:=�o7���a08<��?������N  ��\�S)*5��v�c��L�Q(�z�N���p��V�E"1,�{=�o��m6;��s���G#��R���A��X�f��d����M��y<>?�O'	��Q(4����o��m��}>��o7������Z��q�|��w;�N  ����G��h�j��E"1��[��K�R	�q8��_�����].7�F�A �x��{=�o�����m6��n��b�d����M���|��w;�g�Y���������m6;�����������x�n��e�y<>?�O'��d�i4:=/�K%�i4�}>?��`(����W+��r�s�\��s9����~���s9��W+����l��u:=���{=��w�]�w�].7��q�|/�K��I$�y<>?�G��h��U��z�N���P$29�w;��s��N�����D��H"����C!(�z�g���V�B��P$��|��w;�S�T
%)��U�u�����w;�S)�j
�R���A ��\��s�\��i4:��O'��B���H��Q�t-+����Q�t-��u:�^�����\�S)*����S)�j�e����O�S)��U*�Z���x�����_�W+��E��x�n�E�q8<>���w;'��d�i�z�N�C!����E�q��^��c1,6��n���Q(�z�N�A��X�f�I$29�w;�N�C�P$��|�o���v�M�s�\'�I�r�f	����T�e2���G��h*����S��J!(��]�w��n�K���d)������U*�Z��q8<����o7�F���P$���^���p�l�k�Z���x��W��j�J���`����f	����T����l�k5�m6;�g�����e2�\���y��_���u:=/�E"1,6�]��{�^������N�C���D!��T�e�y���o�[-+������T
%���E"1��V������D����L��h��U*5-�k�������Z��C!�h��z�S)�j�e�y<>�_/��e29�n���r&3�L���x�w��n��e29�n��e29.�[�V��b�H��x�w;�����^��a��\�g3�������L#�H��Q(4:���g3�f�D���X&3&3�s9��{=�W+�J�P����d�i���n�K%)���]��{���g3�L#$29�w��n�K%�i4�}>?�C�P�d��J��p,6;�S)*5��v���a�x���k���f��d��J�B ��X&3���C��H�b$29��{=�o�[�V�a0���O'�D!(��]�����_�W��j
%�i4�����w;��G��h�u:��O'���R	"1,6�].7��f	�b����A 08��_/!��T�e2�\�S�T
��I$2��N�`�h���j�J�a���N�C�P$29.7��C�P$�y��_���u:=/�E"1���K����������R	�q�|��k�����i�z��G#����d)�j�J���`(�z��G��h����n�B�`(4�������}�?�O�S�T�e��|/���Q�t����m6;'�I$2��N�A���L�c�X�s9�����z�N��a�x.�[��K%��t���[-��u�}�����o7���a��\�g�Y,6�].�[-+�e��|��w;�g�Y,6��n�E"��L�������c1�v�Q�t�m�{�^�G����J�a���N���P����V����h*�Z�Q����f����I$29�w�].��������m6;���y�~�O��i4:���g���V��b�H"�X����t�m�{=/����Y�v��C�P$2����c�X�s�\�����^�G#��R���A�p,6���W�U���].7�Q(4:=�o7�F��`��Z�F  ��\��s�\�����^��`����E����N�C!���J��A�p�l���z�N  �x���k5�m6���W+��E�q8��_/��e29������o7�M�s9.�[���e29��W�U*5�V���Q(�z�N��a��\'��d)������U�u:��O'�������D�a0�|��w;'�I��������Y��[-�k�Z������b�H"1�v��h*5-�k�Z�F  ������q���O'��B�@  08�~���s9�����z����q8��_/��A���L��h�j��r�L�Q��Z��h��z'	"1,�{=��k����S)���j�e29�n�K%���Z�Q(4�}���o7�F��`�t�m����_���u��~��g3����a0��^ ����F���P$2�\��s9�n�K�R��B�`��T
��I$���^�G#���B�`(�����k�Z�c1,6;�g3�L��q�|�o��������m6�].�[���e29�n���r��S�T
�R	�q8<����?�O�S)��U*5����m�{�^�C!��Z#���I����V�P�d)�u:�^�G�Q����f��d��J�B��P����d�i���n��e29���k5����m6��n�E��x��{��O'	"1,��}>?��a�x�n!�t����m��}>��������o7�M&3�L#�H�b�H�q8�~�O�S�T�e��|/�����T�e���^��c1���m6�]���}��_/���r���i4:�^��c��L�c�����a�x�n�K�R��B�`�h*5�m6��n�K���d�i4��~��g��l+�e�y<>�_/��e��|����}�������?����x����~���s9��{�^��P$2�\���y�~��a�x�����_/�E"��L���T���Y,�����o7�M&3�L�c��L���T�e�y<�?��c�X���i4�}������o7�F���@��P��R��B�@�`(4:=��k5��v�M�s9�n��A�p��[-�U*5�m6����������k5��v�F�@ ��X��S)*5��v�F���H��Q(4:��O'��B��@  0��^��c1��[-���z��G�Q(4�}>��o7�c�X���i4:��O'�����d��t-�U���]�w;����q�|�W+�J!��T
���d)�j��E�q8<�����o7�F  0�����s��N�@�`�t���[���e�y<�������?�G�Q(4�}���_��k5-�U*��M�������s9�n��e2�\�S)�����j��r��y<>����{=�W�U�u�}��?�O'��d�i4:=�o�[�V�a08��_��k5��v#$��|����}�?�G�Q(4�}�����?�O�S)�j��r�f��B���@�`�t�V�E"1�l��u:�^��c1�l+�e29�w��n�K%�T
%)���j�J�B���@  08�~�A�p�l�k�Z��C�P�d���Z�F��`����E"�X�f����`���J���`����f�D�a08<�?�G#$�����g��l����]���}>��o�[-��j�e2�\��i4�}�����{=/�E"1,6;��G�Q(�z������\'��d���Z�c1�l��u:=�o7���T
%��t-+
%�i�z'��B  �x���}>��o7��f	����N��`�h��z��G�Q(4:=���{=��k���f�I$��|���{=���{=�W���U*��M&3������X&�Y,6;�g3��F �p�l������j��E"����C!�t��K�R	��������Q���M��y��_/�K�R	�b��D!��T
%�i�z��G#�H��Q(4:=�����~�G�Q���M����^����X���i��].�[-�U�u�}�?�C��H������c����C!(�z�N�@�`�t�m�{��O�S���E�q8<�?�O'�D�a�����c��L����\���y<�?���s�\�S)�j��E"1����v��f���R��B ���L�c1��[�V��������A �x��W+�J���`�t��v��f�I�r�L�Q���M&3�L�c�X�f�I$2�����q��^�G��h*��M&3&3���i4�}>�_�W�U*5-��u��~���s9.�[����r�L���x�w;���c1���K%)��z�N���p�l��u:��O�S�T
%)�j
���d�����f	�b�H"1���m��}>?�C!��T�e���^��������P�d����M&3�L��q�|�o7�M&�Y����v�F����@�`(4�}>?��`�t�V��b�H�q8<>?��`�h����U*��M��y�~�G#�H"1�v�F����@���H�q8�~���p,��}>?��g�Y,6;�����x�n������J����P$2�\������O'�I���l+�J�B�`��Z��q���O��i��]������o7���a08��_/!��T
�R�D�a�x�w�]��{���g���V!�t��K%��J!�h��z�g��l�k5�m6;���c1�v�F�A 0�|�o7����i4�}>?��g3&���V�E�q���O'��d���Z�F��@  ��\��s��N�C!�����b�H"1����e2��N��a08<����?�@����D�a0��^�A���L#�d��J�B ���L�c1��[��K%)�������u��~�O'�I�������r�f	���h�u�}>?��c1�l��u:=���{�^����X&3�����O'	����T
��I$�y���o7����J�B ��X�f	���\'�I��������Y�v�����t-+�J�P���I$��|�o�����m������w��n���r�f�I��Y�v�M&���V������C��H�q8<�?��c�X�f��d�i���n��e�y������}>?��g3��F����@��P���I�r�L#�H"1�v��f�����d)*��M&�Y,�{��O�S���E�q��������^�G���T�e2�\�S)�u:���g�Y,6�]����~���s����c1�l����]��{=/�K%���Z�Q����f��B���@  ���N��P�r�f����I��Y��[-�k�Z��C�P�r�L�c1��[�V�E"���F�A 0�|/���`��T
%��t-+�e29.7��f�I$���^��c�X�s9��{=�o7��f��d�i�z�g��l�k5�V���X�s9.7�F�@�`(��].�[�V����P$29�w;�N������F�@�`�t���e�y<>���w;�N�C��H��Q(4:=���{=�o7�����t�����v�����X��y<>�_��k�Z�F�`�h���j���Y��[�V�a��\�g�Y,��}����o��m6;��i�z�g��l+���b��D!(�z�N��a����G�Q(����W�U*5�����v�M����^��c1�l�k5�����v�F��`�h�����W+���Y�v��f	��Q����f	"1�v�M����^���@ ��X���i�z��G�����E"1,�{=�o7��q�|�W�U�u:��O���t�V�B�@�`���J�����H"��L�c���F�A���L#���B�@  08<>����{=�W�U*�Z�F�A 0�|�W+��E��x�n�K�R	�q�|�o�[-�U*5�m���~�O'��B�@  08<����_�W����j��E��x�n��e�y<�?��`��T
�R����`��T
�R	�b$��|������_/�K��I�r��S)��z������O'	���h*�Z�c���F�A�p�v��C!������Q(��].���v���S)����U*5�m6;�N��a�x��{=����z��s9�w;'�D�P��Y�v��C!��Z���a��\'�I��Y,6����k���f�I�r���i�z�����x�n�K���d)�j����l+�e29������o7�F�A��X�s9���k5-�k5��v���a08�~�G#�H��Q�t�m6��n���`�������h�u�}>?���q8<>��o7�M��y�~��a08<>����{=�o�[��K%)*�Z�c�X&3��F �p�v�F��`���J��A 0��^�`�h*�Z�F��`(�z������\'�I��Y,6;��i4���_/�B�@ �p���m��}�?���q����g��l����].7��f��B���H�b�H"1,6;�N�C������`(�z�N��a08<>�_/�E"���F��`�h����n�K%��t��v�F�A�p��V���Q�t�m6�]��{=/!�t���[-+����Q�t-+�e29�n�E"��L�Q�t��v���S)*���f���R	�q�|�o�[�V����h��U*���f��d)*�Z�c1,���~�C!�h����U����n�K%����b�H"1�l��j�J�B���@  �x�n���r��S�T
%)�j����Q�t�m����_�W�����U������k5�m�{�^��c���F��`�h�������j�e29.��m��}�?�G#�r��F�A����F��P��R�D�a0�����s��N��`��T
��I�r�f����`�h�u:��O�S)�u:���g�����e2�\�S)�j��r�s9����~�����|/�����T
�R	"1���K�R	�b�H�q���O�����M&��l�k�Z�c1,�{�^���p�l��j
%��t��v�M��y�~�O����Z�F��`�t�m�{=/�E"����C!���J�B  08�~�O'��d)*5�m�{=/�K������d�T�e29.�[-�k5���[-��������u��~��g3�L�Q(��]�w;�g�Y,�{�^��a�x�����_�������W������j���Y,��}>?���s������x�n����Y�����[-+���b��D�P�r�s9�n�K%�i�z�N��@��P��R��B �p��[-+��r��S)�u:���g�Y�v���T
%�i4:=���{=�o���������v��C!�h�j
�����I���l+�J�a�x����u�}��?�O'	"1,6�]��{=��w;�N�C!(�z'��d����M&3�L�c�X�s�\�S�T
���d)��U�u:�^�G���T
%�i�����k�Z������L�c1�v��f�D���X�f�������I$�y��_��k5���[-��u�}���o���v��q��^�����\��s��N�A������a0���O'�I$��|����}>?����X�f�I$�y<����_�W�U����n������D�������a���N�A �x.7���S�T
�����I$�y<>?�C��H�q8��_�W�U�u��~�����\��i�z�N��@  08<>?�O'�I����V�B��@�`�h�j�J��p,6;��G#�H��Q(4��~�G��������h�j�e29�w;�N �����C�P��R���A 0�|/������V�E�����G������b�r&3�L���x.���v#��R���A 0���O�S)�j
����R��B  ��\��s9�n��H�b$�y��_/��H�b$29�n�E��x��W+�J�B �p��V��b��R�D!��T
%�T
��I�r�s�\��s9�w;�N�C!�h��U*5-+��r&3�f	�q8���o7���S)�u�}����?�������O'�I��Y,�{=��w����k�Z�������c1��V����L�c1���K����R	��Q(4:=��w�]�w�����u:=��w;'��B  �x�n�K��I��Y�v��h�j��E"�X��y<��?�O'��B�@  �x�n�K%��t��v�M&����K�R���A�p�v����p�l+�e2�\�g�Y�v�M&3��F��@��P��Y�v��C�����A �x.7�M�������s�\���y<��_�W+�e2�\���t���[-����].7�M�s��N���p�l�k5��v�M�s9.�[����r�f�I����V�E�q8<��������o��m6;�N�C!��T�e29.��m��}>?�O'���A����F�@�`�t-+�J��A 08�~�O'�D��p��[-���z'�D��p��V�E"��L�c���F �p�����r���|/�B��@  0�|���{���g��l��u�}��?�O'	�b�H�b�r&3�L�Q(�z��s9�n��b��D�a0���O��i4��~����H�q8<>�_�W�U�u:=/��A�p�l+��E"1��V��b�H�b��D!���J�B�����B �����C����B�@ �p���K%��J��H"��L��q8<��_/��e�y<>?��������`��T
�R	�����J�B��@�`(�z�N�C���D���X�f	��Q���M&����K�R	"���F��`(�z�S)��U���]�w;���c�X��S)��U���]�w;�N�C��H�b���l�k�Z���a08<>?��g�Y����v��f���R	�b���������I$�����g�Y,�{�^�A�p�l�U�u�}>��o7��f�D����L#�H��x.7�c���F�@�`(4:=�o7�M&�Y�v��C!��T
���d)�j�e�y<>?���s�\�S�T���Y����v�M�s��N  0�|�o7������L#$2�\�g��l�U��z������O'�I�����K%�T��r�f�I$��|�o7�M&�Y��[-�U�u:=/�B ����F  ��\�g��l��j�e2��N����X&������r��F�A��X��y<>?���s��N�C!(�z���y�~�O�S)�j�J����P�d)��U*5�V�B��@  �x��{�^��`���J�B�@�`(4���_��k�Z�c1��[-��j
��I$29.7�M�s�\'�I�r����a��\����Z�F�A �x.7���S����b�d�T
%�i�z��G����J!���M���|���u:����s9.�[�V�B�`(4���_��k5��v�F���@  �x��{�^�G#�H����T�e2�\�g3��F��`(�z����q8<��?��c�X&���V�E�q8�~ �����C!(�z���y<>��o���v�M&�Y��[-��u�}>��o7#�H�b�H"1�l�k5����m�{=�o7������L#$2��N���p��V�B�����@ ��X�f�D��p����e29�n�a�x�n��e���^�G��h�j���b�d���Z������G#���B  ��\'	�q8�~�G#�H�q8<>?�G#�H�b��Y,6;�N���P��R	�q8��_/�K��I�r��S�T���Y���m��}�����?�O�S��J�B���@ �p�l��j�J��A�p���K��I$29�n�E"�X��y<�?�O�S��J����B �p�l��u�}�?�`(����W+�J���`(�z���y<��?�O'��d��t��K���d�i4:=�o7�M���|���{��O'�D������`�h���].�[�V�E�q8�~�O�S)���]���}����?�O�����M&�Y�v��f���A��X�f��d)�j�J���`�t-��j�J�a�x.�[-+��E"1��V����h��U������k��M�����O'�D�P�d�����f��B����@ ��X&3&3�L#�H�q�|�o7����i4:=���{=����}>����{����s��N����X��y<>?���s9.�[����r�����p�l+�J�B  08<���?�O����Z��q��^�G�Q(4���_��k5�m��}�?�O�S������h*���f�I�r��F  �x��W+���������b�d��t�V��b�d�i��]��{=�W����j��E��x��W+��r��F�A��X&���V!(�z�N���@  �x.7���S�T
%�i4:�^�@  �x��{=�W+��E�q8�~�`(��]�w���W��j
%�T
��I��Y,6��n��b�H�b�d)�j��E"���F��`���M�s�\'	��Q��Z��C!���J��p������Y�v������L�Q��Z��h*5��v�M��y��_/�K%�����Q��Z�c1,�{=/�K�R��B��@ �p�l�k5-+�e2���G�Q(4:���g��l�����n�K�R	�b�H���\���t�m���~��a�x�n�E�������q����g3�����O'�I$29�����_�W+�e�y��_�W+���Y�v�M�s����c��L#�d��t��v�M�s�\�g3�s9�w����k�Z�������F��`�t�����v��q�|/�K%��t�m6;��G�Q(4:�^����x�w;���c1�l�k5-��u:=����}>�_/�K%�T�e29.7�F�A�p,6�����u:��O���t��v�M�s9�n���r�f�I�r�L���x�n����h�j�J�a�x�n��e��|/�E�q8<��?���q�|/�P�����R�D!������i4:=�o��m��}�����������o�[-���z�g���V��H����N�����L�c1��V����P$��|�o����[��������K�R	"��L#��D�P�d�T
%)�u�����w�].��m�{=��k�Z�������F���H�b��R���A 08<���?�O'�I$�y�~������^����x�����z�����x�n��b��D���X�f���R�D!�t-+
�R�������D�a�x�w;����q�����s��N�C�P��R	��Q(�z�������S)*�Z�c�X�s9�n��e2�\��i�z�N  08�~�G#�H��x.�[�V���Q�t�m���~��g3�L�c1�v��C�P��Y��[�V�E��x.�[-+
%�i���n�a0�|�o�[-+�J��A ���N�A����F�`�t�m6;�N  08�~��c�X�f��B�����@�`�t-�k���f��d)�j��r�L#�H��Q(4��~��g�Y,6�]���}>?����x�n�E"���F��`��Z#�H��Q���M��y����w;�S)�u:=��k������t�m6��n�E"1���K�R��B��@  08�~�O'��B�@���H"�X&3������X&3���C�P$2���G�Q(4:�^�G#$29��W��j
�R	��Q�t�V��b�r��F�@ �p,6���W+
%��t-�k5��v�M&3���C��H��x���k�Z�F��@����D�a���N���p����e2�\�g�Y�v��f���R	�b�H����T
�R	�b��R�D�a�x�n�K��I�r��S��J�P�r��F��@���H"�����a08���o7�F�`�h��z��G#�����R�D��p��[���e29.7�c���F�A�p��[�V�B����@��P�r�f�I$2�\���t�����v��f�D�a��\'���R�D��H"1,���~�����|��w��n��e2��N�C�P��R	"�X&��l+��r��S)��U�u:=/��e2�\'�D!�t�m6�]���}>��o7��f�I�r�s9.�[-����j���Y,����_�W������j�e2���G#�H"��������L#��D�P��Y,6�]��{�^��`(�����k�Z�Q����f�D�a�����c1��V�B�`��Z�F��P�d�T
��I$2���G�Q�t�m��}>?�G#�d)�j��r��S��J�B�@ �p��V���`(4:=���u�}����w�].�[��K%��t-���z'��d�i4:=���{=��w��n�K%�i�z���c1�l�k5������[-�U��z�N�C�P���I�r�s9�n�K%�i��].7�F�`�t��v���S�T��r�L�Q(4�}���������o������v�F�@�`���J�B���H�q�|�W+
��I��Y,��}�?�C!�h��U*5�m�{=�o���v�M&�Y,���~��g3�L�c�X&3�����p�v�M���|/��p�l+���������Y��[�V��A 08�~�G#�H�q8<>�_��k5��K��I��Y,6;�N��P�d)��U�u�}>?�G#$29��W�U��z����|�W+
��I$��|�o�[��K%�T
%��J!��T��r�L��q8�~��g3�L�����E�q8��_/�E"1����e�y<>?��g���V�E�q8�~��c�X���i4��~����y<��?�O'	�q��^��c�X�����O��i�����k�Z��q8<��_/�K�R	�q8�~�C!�h��U�u����o7��f�D!(4:��O'��B�`�h��U*5�m�{=����}������{=��w;�N��������`(�z�N�A 08<>�_/�E�q8<>�_����z�g3&�Y,�{=��w�]��{���g3���C�P���l�U*5����r��F�A�p�l+�J��A����F�@�`��Z��C�P��Y�v�Q(4:=�o7��f	"�����a0����g���V!��T
�R�D���D��p�l���z�N�A�p��V���`�h�j�J�����H��x��W+�J!(4�}>�_�W�U*5�m6;���t���������[-+����Q(��].�[�V�E�q�|�W+�J�a0�|/��b�H�b�H���h*�Z�����N�A�p�l+��E�q��^�`�t��K���d)*�Z���x�n�P���l����].�[��K��I�r�f�D��H�q���O�S)���]���}>���w;�g��l�k5�m����_/�a0�����s9�n��e2�\'�I���l+�e29�w�].�[�V��b�H"1�v�M&3�f��d�i�z���c1,���~���q8��_/������J�B�@�`�t��v��f��d)�u:���g3��y<>�_/���r�f���R	"1,6;�N�`(������u:�^��`�h*5-��u�}>�_/�B  �x����������u���_/�E"��L����\'�D�P$�y�����{=�����~�O���t-���z�g�Y�v�M�s�\����|��w��n�a����G�Q�t-+���b��R	"����C!��Z�F�@  �x.���v�F���P$�y<����_�W�U*5�V���`�t���e2���G#���I$29.7���x�w;��G�Q�t��v�F�@�`��T
��I$�y<>?����������y�~��g����K%��J��A�p�l�U�u��~���s9.��m6�]�w����k5-�k���f���R�D�a0��^���p�l�U�u������{=�������W�U*�Z���a08�~�O�S��J���`(��]�w��n�E"1�l�k5-��j���b��D!(4:=/������V��p��[-��������u:=/���r�s9.�[��K�R	���\�g�Y��[�V��b�����`��T�e29.�[-�k��M�s�\'�����P���I$�y<�?�����|�W+�J�P�r�f	�q����g�Y�v#��D�a0�|/�K�R	���h�u��~�O��i4�}>���w��n��p���K�R	��Q(���n�K���d�i��].����[-���z���c�X���i�z��i���n�K�R��B �p��[-�k�Z���a�x�n���r���C�P�r�L����\'���R��B�@  0��^ �p���K��I�r�����Z#�H�q���O��i�z�g�Y��[-�U*5�m�{=��k5-�U��z�N�C!��T
�R	�q��^������A 0�|��w;���c1�l�U���].�����m6������z�g����K%�����f���R	�b��D���X&��l�k5��K�R	"1�l+��E"��L���x�w����k5�m6;�N  ��\��s��N��`�t�m�{=�W��j��E�����G#��R	"1,������w;����q��^�A�p�l����]��{���g�Y,�{��O�S��������J����L#$��|����z�������N��@�`���J���`��T�e2��N��a�x�����z�S����b�����R	�b���I$�y��������_/�B�����@ ��X&�����e��|����}>�_/���r����t���[�V��b�����R	�������q8���o7�M&�Y�v�M&3���C�P��R����`�h��z�N�@ ������a0�|�W�U���].7�F�A�p,�{�^��a08��_/����Y����v�F�A���L�c�X��y<>��o��m�{�^��������@��P��R�D���X�f	���h��U*�Z#��R������H��x�n�B��@  ���N��a0���O�S)����U*����S)��U��z��G#$2�����q�|�W+
%�i4�}����_/�K%�i4:=/��A 08�~��g3��F�A 0��^�G#�r�L�c1�l+�e2�\�g3��F��`��Z���T
%��t�m6�].7�M����^�A����F����H�b����A 0�|��k5��K%���Z�Q�t�m6;�S�T
%�i4�����w��n�K%�i4�}>��o7��C�P�������d)��U��z��s9.�[-���z�N�A��X�f����I$���^�@  08�~�G�Q�t�m6�].7�M&�Y,��}>?��g�Y,�{��O�S)��U�u:=�o7�F��`(����W+
��I�r�L#�H��x�����z�g3��S)��U�u��~�G#�H"��L#$29�n�E"�X����t��v�F�`�t��K%�T����l�U*�Z�c�X��y<��?�G���T�e�����g3�L��q��^����H��x�����z�g�Y�v�M&3�L�Q(��].7�F  ���N������F�A���L�c1�l��u:�^��a0�|�o7�c��L���x�n��e29�n���r&��l�U*�Z����p,�{=��w;�g3���C!��T�e29.���v�M&3&3��S����b��D��H�b��D�a�x�n��e2���G�Q(4:=��k5����m6;'	"��L#����A ���N�A ����G�Q(��].7���x�n�K�R	�b��D����L����\'�I$29�����_/�K��I$�������y�~�G#$�y<>����{��O'���R	����T��r����a�x��{=���{=��w�������].�[-+�e�y�~��g3���C���D������C�P��Y��[�V�E"1�v�M&3��y<>?��g3�L�c1,6;�N��a0���O'��d�i4:=�o7�����X&��l��u:�^�G#��D�a��\'	"�X�f	����T
�R�D�P����V������J����P�d���Z�F�@  08�~�G��h��U*5�m6;���c1�v������Z#�H"���F���@  08<�?��a������q8<�����w;�N�A��X�����Z����p�l�k5�V��b$2�\�g���V���Q�t�m���~�G#�H�b�H��Q���������M&3��F�@�`�h*��M&3�L#��R�D�P�r������M&��l�U��z��G#��Y�v����i�z�N�A�p,��}�?����y�~�A ��\�g3��S����b�H��x�n��A �x��{=��k5-��j�J��A 08��_/��e��|�W�U*��M&3��S)��z�������g�Y,�{���g��l���z�S��J!��T
�R�D!(4�}>�_��k5��v��C!�h*����S����b�d�i�z'�����P�r��F�����D!��T
��I$�y<����o�[-�k5-����].��m6��n��e�y�~�O'��d����b�H�b$2�\�g�Y��[�V�����H"1�l+�J!���J��p��V�B��@ �p�v��C!�h*��M&3�f�I$29�n�E�q8<�����{=�o��m���~��g�Y,6������z�g��l�U�u:�^�G#�r��S��J���`(����W�U*5��v���S��J�����H��x�n��b��D��p,6;�N���P�d�i����W�U�u:�^�G��h����U*��M&�Y�v��f����I$2�\�g�Y,6;�g�Y,6�].7�M�s����c1,�����������o���v��q8�~����y<��?�C���D�P�r�L�Q(4:=/��b$29����u�}��_/�K��I��Y��[��K%��t-�U*5-�U�u:��O'�I$2�\���y�~�O��i4�}�?�@ ����F�A 0����g��l�U����n�B  08<��?�G����J���X&�Y��[-�k��M&3�f�D!�h*5��v�F�A �x.7�F�A���L�c1�l�U*5-�U*��M������g3��S)��U�u��~���q��^�G#�H"1���K%���Z����p,6���W+����Q(�z����Z�F��P��Y,��}>?����x���}>?�O��i4�}�?���q�|�o7�F�A�p�l�U*5����r������X�����Z#���B�@����D!����f��d)�u�}��_/�E�q�|�W���U��z��G#�H"1����������v���a��\'��B��@  �x�n�K��I�r&�Y�v��f�D�a�x�n��e�y<>�_/��p�v�Q�t-�U*�Z#�����K��I$2�\��s��N��a0��^�@ �p���K%�T���Y�v�F ������a08<���o�[�V�B�@�`����E"1��[���e29��{��O'	�q8<>�_/�K�R�D����B���@���H"1��V�B�@  0�|�W+�e��|����z�g3�f�I��Y,6;��s���G�Q�t�V���Q(4:=��w�]�w�].7��q8<�?��g3�L���x.7�Q������i4:���g3�L#��D�a0���O'�D�a08<����w;��s�\'�I���l+���Y�v�M�s��N����X��S)*5��K��I$29���k��M&�Y���m6�].7���a08����w�].7�M��y���o�[�V��A������a��\�������S�T�e2�\�g��l�k�Z�F�A��X�f	"�X�s9�w;�g�Y,6�].�[-��u:=������n��b��D�a��\��s�\�S)�����j�J�B  ���N�C��H���\��s�\��s���G�Q�t-�U��z�N�C!(���n��p�v���S)��U*5�m�{��O��i4:���g3&����K��I$�y���o7�F �p�l�k�Z�Q�t�m6�].7�Q�t�����v�M��y<�?�G#�H"1��V�B�@ �p,6��n����Y,6�]�w�]���}>?���s�\��s9��W+
�R	"�X���i��]�w;�g�Y��[-�����n�B����@����D�P$��|��k�����i4:=/�E�q��^�C�P�d�i��].��m6��n�E"1����e29.7�M&3����t�V���`��Z�F���P�d)�j�J�a�x.7��f�I��Y��[-�k��M&���V�E"1�v��f���R��B�@  0�|��w;�N��@��P�r�f����`��������Z�F�@  ���N�������A���L�Q(�z����q8������}>?�O�S)��U*�Z�F ��X&3�L�c���F�A �x�w�]���}�?�G#�H"1�v��C��H��x.7��f��B��@  0�|�o���v�����N�������C!�t��K�R�D��p�l���z��s�\�g��l+�e��|���{�������^�G#�H�q8�~�A�p,�{=�W+������T�e2���G�Q�t-���U����n�E�q8�~��c1����e29�w�].7���S)�j��r�L���T�e��|��w;'���A ������q��^�C!��T
�R	"1����e29�n����Y,6�].��m�{�^�G#�H��Q(4��~������^��c1��V����P$2���G#�H�q�|�o�[-���U*��M&3�L�c�X&���V�E"1���K%��J�P$29�w����k���f	���h�j�e29�n�E�q��^�G��h�u�}�����?����x�w�].7�F�A�p�l+
�R	"1��V�B �p,6��n�B�@�`�����b�r��S)*�Z�F�A�p,6;�����^���������p,6;����q����g3�L#�r&��l���z�����x�n���r���C�P���I��Y,�{=��k5���[���e��|�o���v���x�n�K��I$2���G��h�j��r&����K�����I��Y�v��C����B�`��Z���T
%)�j�J!(���n�K����R�D�a0��^�C!(�z������\�g3�f�I�r�s��N�C!��Z�c1��[-�k�Z���x.��m6���W���U*��M�s�\'��d�i��].�[�V�B�`�t�m��}>����{�^�G�Q(4���_/�K%�i���n�����H�b�d�����Q�t-���z�N�A�p�v�M&3&�����e29������].7������L#�H�q���O��i4����o��m6�].�[��K%���E"��L��q��^�A 0���O'��B��@�`�h*5�m�{=�W�U*5����m6�]����~����y<�?����y��_/�K%�i�z�S�T
%��J����L���x�w;'���R�D!��T����l�U��������z������f�I�����K���d���Z�Q��Z�F�������A���L��q�|�o7��C���D��p�v���a�x�n�K��I$2�\'�I��������Y,���~�O'������H�b$�y<����o7��q8<�?����y<>?�������@����D!(���n�E�q8�~�`�t�m6;�S)*��M�s9.7�M&3�L�����N�C!����E�q8�~�O'������H"1,��}�?�O'	��Q��Z�F�@  �x�n���Q(4��~���p��V�E�q��^����x������].7�M�s9�w�].�[�V!��T�e29���k5����m�{=���{=��w;�N  08<���_�W+��E"1,6�].7����i���n�K%�i4�}>?��g3&�Y�v#�d)*��M&3��y�~��g3����^����X���i�z��G�����E"�X�f�I$29��W�U*5�m6;��G#���I$��|����}�������w�].�[���e29.��m6�]�������w;�g3&���V�����T�e�y�����{=��w�].�[�V!�h���j����Q��Z#�r��S���E"�X�f��d����b�����K����������R	���\��i4�}>�_�W+��r�����p����e29.7���a08��_��k��M���|/�E�q�|�o��m�{=/�K%�i���������n�K�R	�b�r����a��\�����M&3��F�@  0�|�W����j�J�B��P��Y,6;��s9���}�?���s9���k�Z�F  0����g3�L�Q��Z���a0���O���t���[-�U*5��v�F�A����F�`����E�q8�~�O���t��K%�i�z'	"�X���|�o7���S)*5�V�E"1,���~��`(4�}��?��c1�l����j��E"�X�s9��W���U���].7��C�P$����O'���A��X�f��B�@ �p����e29�w;��G�Q�t�����Y����v�M���|/�E�q�|��w;�g�Y,�{=/���r��F��P������e29�n���Q���M&�Y,6�].�[-+���������b�H��x�w�].7�����E"1,��}>?�C!�h��U*�Z#��Y����v����i��].7��C!���M&��l�k5��v�M��y<>���w;�N�`�t�m6�]��{=��w;�N�A 08<>��o�[�V�E�q8<��_�W�U�����W��j�J�B  0�|�o7�F���P��R�D�P��Y,��}���_�W+�J�B��@  0�|��k5�m�{�^�@��������P$��|/����P��Y,��}>������~�G��h���j����Q�t�m�{�^��a08�~�O'	�b����A��X&3������M&�Y,6������z�N�C�P�d�i�z�S����b��D�a�x��W��j�J�B���H����T
%��t�V�B��@���H���h*5-���z�g��l����j�J�a�������x�n��b��D!�h�u:�^�C�P��Y,6�����u:�^��c�X&3��S)*5�V�B�`�h��U����n���Q(4��~����x�n�P�d�i4:�^�C!�t���e�y�~���s9.7�F �����C!(�z�N  08<>�����}>?��c�X��S)�j
��I���l�U*5-�k�Z����p�l����].���������v�F ����F�������@  �x.�[�V�B������A ���������N�A�p��V���X&�Y�v��f�I$�y��_��k��M��y<�������o7�M&3��F�A �x�n��e�y���o7�F��P�d�i4:��O��i4��~�G�Q��Z�c1,��}>����{�^���q��^�G��h�j�J�B���@ ��X&3�L��q8<>?�G��h*5��v��f	���h*�Z#��D!��Z��C!��T
�R��B �p�l�U�u�}>?��@����D�P��Y,6��n!�h�j
%)�j�J��A��X�s9�n���r��y<>?��g3���C�P$�y�~���q8<��?�����|/��e29.7���a�x.7�F��@  �x.���v�M&3�s9.��m���~�O'�I�r�f	"����C!�h�u:=���{=�W�U��z�N��`�t�V���Q���M&3�f��d��t��v�M&��l�U*5�V�E�q8�~�O'	��x.7�F�����@  0����g�����e������s��N��@  08<����?�@�����B��P$29.7�F�A���L#�d����M&����K%���Z�F���������P�r��S)�j��E"�X�f��d)�j�J���`���M&3��S�����Q��Z�F�A�p,6������z��G#�d�T�e2����c�X���i4�}>�_�W+��E"1��V���������`��Z�F���P�r�f��d)�j
��I�r�L��q8��_/�B�@�`(4���_/����Y���m6����k5��v�M���|�o���v�M&3���i�z�g3��F�A�p�l�U*5��v���S�T
��I�r�s�\���y<���?���q8����w���W�������U����n���r�f����I$��|�W+
��������I$��|����z���y<����_�W��j��E"�X&�������Y��[��K�����I$���^���p���m��}��?��g3�L�c1�v��f����`���J��A����F��`�h�u�}�?�C!�����b$�y���o7������Z�F����H��Q�t-�U*���f	"1�v��f�I���l�U�u�}>?�O'��d�i4:=�o�[����r��S����b�H�q8�~����@��P$�y<>?�O'	���\���y�~�G#�r�����Z��q�|/�K%)���j���b��D��H�q��^�G#�d��J��p,��}>?��c�X���i�z�N��a�����c�X&�Y�v������L��h�����j
%)�j�J����B�@  08<����w�].7�M�s��N�A�p�l�k5-�U�u:=��k5��v�M&��l�k�Z�����N��`(4�}�������w�].7�F��`(4:=��w;��G#��D�a0��^��a0����g�Y,������w;��G�Q(���n�E"�X&3��S�T
�R��B �p��[-��u:���g3�f��B�`�t������l�U��z����|��w��n�K%�i�z�g�Y��[-���U��z���y�~�O'�I$�y��_/�E����N��a08���o7�M�s��N�C�P$��|��w;����|/��e��|��w;��s9��W�U�u:��O��i4:�^�G�Q(4:=/���r&3�L�c1�l�k���f��d���Z�F�A �x��{=��w������z�N��`(4:�^�G�Q(4��~��g3�f������R	"1��[�V��b$��|�W+�J�a0��^����X&��l��j�J�B�@��P$�y<>�_/��e2����c1,6�].7���S�T
%)��U��z��G#���I�r�L#�H��x.�[�����Y�v��C��������H��x.����[-�k�Z��C!��T
������d�i4:�^��c1�v�F�@ ��X&3�L#��D�P$29���k��M&3�s�\���y<���?����x.7�M��y�~��g3�L#�r��F  ��\���y<>�_/��p��V�a08�������~�O'�D��p�v�F����@  ��\�S)*��M&�Y�����[-�U��z��G#$�y<>?�G�Q����f�I�r��S�T�e2���G�Q�t�V�����T
�R��B ���L#�r�f	�b�����`�h�����j�J�a����G#�H��x.7�M�s9�n����P$�y�~�G#���B  ���N�A 08�~�O'	���h*5-�U��z�����x.�[-�k5-���z�g�Y�v�F�A�p�l�U�u�}>?�����|�W�U�u:�^�C�P�d��t��v��q8<��?��g�Y���m6;�����^����x����u��������~�O�S�T
%�i��].��m�{��O�S)*5�m6�]�w;�N�@  �x��W��j��E"1�v�M&3�f	"1�v�c1�l+��r����a08<��_�W�U*�Z��C!(��]�w�].�[-��u:�����y�~��`�h���j���b���l�U��z����|��w��n�E"1�l����j
����R	"��L��q8�~�O��i4:�^�@��P��Y,���~���s�\����Z#�d)�u:��O�����������M���|�o7��f�I�r�L���x���k5-+��E�q8�~���s�\���y<�?�G��h*5��v��C�P�d)���].7�M�s�\�S��J!�h�j��E�q�|�����~ �p,��}>����{�^����x�n�����l+���Y,6�]����~���@ �p,6;�S)*�Z�F��@ �p�l�k5�m6�].�[��K��I����V�a08����w;���c1�����r���C!�t-�U�u��~�O'��d��J�B�`�t-+����Q(�z�N�C�P�d��t�V���Q�t-��j
%��t-�k5�V��p�����r�L��q8<��?����y<�?�C!��T
����R	�q8�~��c1�l�U*5-�k���f�I$2�\�g��l��j����l��j�J�B�@�`�h�j��E��x�n���X�s9��W�����U�u��~��g����K%�T
%���Z�Q���M&��l��j���Y,�{=��w��n����Y���m6;�S����b�H"1�����r���|�����]�w�]�w�]����~�O'��d)�j
��I$2���G#���I$�y<�?��g3���i�z�N��a�x�w;��i��]�w���W���U*�Z��C�P�d)*5�m6;'�D�������a�x.7����i�z����Z�F�A�p�l�U�u:=��w;��G�Q�t�m�{=/�E�q8�~��c1�v��f	�b��Y,��}�����{=/�E"�X&3&3��S�T
%)���j��E��x.�[-+�J�P��R���A�p�l�k5-�k5-�k��M���|�W���U��z���y�~�O�S�T
��I��Y��[������l�U�u��~�O�S�T�e29.�[-�k�Z��C�P��R�����P�d)*5-��u�����w;���y<�?�O'	"1����e��|����}>�_�W�U�u�}>�_/��b���I$2���G��h*���f�D�P��Y,�{����s9��W+�J�����F��`���J�B��@�`�h�u����o7�F  0�|�o7�Q(4:=��w;�N��`(4���_��k���f	"1�l��j
%�T�e�y<>?��g�Y�v��C�P�r���i��]����~��c1�������l���z�N  ��\'	�b�H"1��V���Q(��]����~�C��H�b�H"����C�P�r&3����a08�~�O'	"1,6;'�I$���^���p����e�y���o��m6;���c1,�{=��k5��v#����A���L#�d���E"�X�����Z�c��L#�d���Z�F��`�����b��D���X�f	���h�u����o7�M&�Y,6;��G#��Y,6;�g3&�Y,�{��O���t��v�M��y<>?��c����C!������Q��Z��C�P��R��B�`(4�}>�_/�K��I����V���`(4�}>?�G#�H�b�H"�X�s9���k5-�k5�m6;���c��L�c�X&���V�E�����G�Q(4�}>�_/�E"�X��y<>?����x��W+��E�q����g3���i4�}�?�G������������b�d�i4:=��w�].�[��K%�i4��~���s9��W+��r���C!(4:���g3��F�A�p�v�F�����@�`���M&3�L�c�X�f	"�X�f����I���l�����n�����l�k��M&3�L����\��s�\'���R�D�������a�x�n���Q(��].7������Z��C�P$�y�~�����|�W+��E"�X������g���V�E"�X��S)��U*5��v#��D!�h�u�}�?�O'�D���X�s�\�S)�u:�^�G��h��U����n�E"�X&��l�U*�Z#��D�a���N�C�������P$2��N���p����e��|�����]�w�].7�M���|������_������n��e29.��m���~��`�h�u:��O'	"�X�f�I�����K�R�D����L������G#$2�\���y��_�W+���b�H�b��D���X&3�f���R��B �p�l+�J�B�@  �x��W+�J�a�����c�X���i4�����w;�N���p���K%�T���Y��[-+��E"1�l+��E"1,��}>���w;�g3���C����B  ��\���y�~���s9�w;��s��N�@���H"1�l�U�����W�U����n!(4:=/�B���@���H"��L��h����U*5�m6;'	"1,����_��k���f���R�D�P�d)��z�g3����a�x�w��n�E"�X�s9��W+
%)�j�e2�\�g��l�k�Z�F�A�p,�{�^���p���m�{�^��a�x�n�K%����b$�y��_��k�����i��]��{�^���P�d���E"�X&3�f��d�������i4:�^�G�Q��Z�F�A ���N��@�`���J�B��P��R	��Q(4:��O�S��J��p�l����]���}��_/��e29�����z��s9��W+����Q�t��v�F�A ���N�A 08�~�O��i��]���}>�_��k5-�k5����m�{�^�C����B  0���O��i4:=�W�U*5�m6��n��b�H�����J���`(4:�^������F ���L�c1�l�k5��K�R	"��L��h�u���_/�E"�����a�x.7��f��d��t-���z�g3�����p��V��H�q8<>��o���v��C!(4����o�[��K%�T
�R���A ����G#�r&3&3&���V��b$�y<>�����������}����_�W+
��I���l����].7�F�A 0�|�W�U���]�w;�S)�j�J!�h�j��E"�X&3�L�c1��V�a0�|/�K%�T�e2�\������O'��d��J��������p,��}>?�O���t�m6;������\�����������^�G�Q�t-+�J��A �x�w;���c�X�f�D!��Z#��Y,6���W+�����h��U���].��m6������z�g3��y<>�_��k5-�����n��p�l+��������E"1�v�F��@���H"1,�{=/����Y,6������z�g3�f	"1��V���Q��Z�F�@  08�~��P$���^�A�p�v��f	�b�����`��T����l���z��i���n��b��D�a0�|�o����[-�k5��v�F  �x���k5���[��K�R	�q8��_�W+�e���^��c����C!����f	����T
�R	�b$29.�[����r�s9.7��h*5�V!���M&�����e29.7������Z#�d���Z�F�@  �x����u�}>?�G�Q(�z�N�C�P�d�i���n��A���L#$2�����q��^����x�n�E"�����a0��^�G�Q(�z��i4�}��?����x.7����i4:=�o�[�V��b$2�\'	"1��[-�U��z'	�b����A 0�|�o��m��}�?�O'�I�r��F�@ ��X�f����I��Y,6�����u�}����_/��e�y<��������{�^��c1����e�y�~�A�p��V���`�h�j����Q(4�}���o7�c1��V!�h�j��r�L�c1,6��n��e�y<��?�A���L#��D�a08�~��g����K%)��U�u:����s�\��i��]��{�^��c1���K�R	"��L�c�X�f���A����F��@ ��X�f��d��t-�U*5�m6�].7���a��\�S�T
%��t�m�{�^�G#�d)��U�u�}>��o7�M&���V�E"�X��S)�j�J���X&�Y�v�c1�v�M���|�o�[�V�����F�@  0�|�W+
%�i���n�K%�T
%��J��A��X&��l��j���b$��|/�K�R	�b�d)��z��i4:=����}>��o��m�����o7�F�A����F�A�p,6;���c�X���|�W�U*���f�I���l���z�g�Y�v��f	"�X���i4:=/�K%��t�m6�]����~���q��^�C!���J��H"1,6�]�w��n���r��F�`��Z��C�P$2�\'�I$29����u:��O'	�q8<���o7�M&�Y�v�c�X&���V���Q(�z��G#�d)���j
%)�j�J��H�q8�~���q�|/����P��R	"1���K�����I$�y<�?��a0�|/�K%�T�e2�\'�I$2���G#�H�b�H��x�n�K%�i�z���t����r���i����W��j
�R��B�`��T
�R�D��p��[-��u�����w;'	��x�n!�t��������v��f��d�i�z���y<��_/��e���^��c1�v�M�s���G#�d�i��].7��f�I$���^��c�X&������r��F�����D!�t�V�B��P$�����g��l��j��r�L#��D��������p����e2����c1����e29.���v�M&3��y<>��o7�M&3��y��_/�K%�i����W+
%)����U�u:����s9��{�^��c1,�{=�o�[-��j�����h��U*�Z#�����R��B �p,�{=/��H���h�u�}>?��g3��S)��U*5�m��}���?�O'�I$2�\'�I$2�\�g�Y,6;'��d�i4�}>�_�W+
%�i�z�N�C!�t�m6��n��e29�n��������e�y��_/�E"��L�c�X&�Y,6�].��m6;�N�C�����A���L�c1�l�k5�m6;�N�A 08<�������{��O���t-�������k�Z��q8<>?��c1��[�V�B��@  ����G#�H�����J����P�d����M�s9���k5�m�{=/�E"���F�A��X������M&3���C�����A����F�`�������h���j������T
%)��U���].�[-+��r�s9��W+�J�a��\'�I$�������y<>�����}>?����y<>�_/�E"����C��H�q8����w��n�E"��L#�H�b��D�a���N�C!�t-+
%���E�q8<>?��`(4:�^��a��\�g3��F���H�b�d�i�z�N�����@���H"1��V���Q�t-��u�}>�_/�E������c��L����J!(���n�E"1���K%��J��H"1�l�k5�V�E"1,�{=�W+��E�q��^�G�Q(4�}�����?�C!������Q�t����r���C�����A �x�w�].7�����X��S)*5�m�{�^�G#����d)�u���������_/�K���d�i4��~��a�x��W+
�R�D��������p�����r&3��S�T
%)�����j��E"�X��y�~�G�Q�t-�k5��K�R	�b������P�d��J!���M&�Y,6�].7������Z#�H��Q(�z'�I���l���z'	�q8<>?��c1��V�E"1��[-���z'��B�`(4��~�O�S��J����P��R	�b�d�T���Y,��}>?��c1,6;��i4:�^�����������\�g�Y��[-������W���U*���f�I$2�\���y�~�O'����`�t�m6;�����x����u��~�`��Z�c1��V����B�`����E"���F�����@ �p,�������{�^�G#$�y<>���w�].7����i4:�^��P�d)�j
���d)�j�J�a08<>?�������O'��B�@  ���N����X&�Y�v�F �p��V���Q�t�m6���W���U*�Z��C�P���I$2���G�Q�t-�U*5��K%�i4����o7��q8���o7�����t-�k5����m�{=�o7�M&��l�k5�V�E"��L�c��L�Q��Z#�H"�X&3���|�W��j
%���E"1���K��I$2��N�C!(4:�����y�~�O�S�T
���d)��z'�I����V��p,6;'����I$�y�~����y�~����y���o�[-���U���].7�M&3�L�Q���M&�Y�v��f�I�r�f�I$2�\'���R	��Q�t�m6�]��{=�o��m��}��������_/���r�L��q�����s9�n��e��|�W�U��z�����x�n�E"�X�f��d�T��r�L#������P��R�D��p��V�a��\'�I$2��N��`(�z'�I$29����u:�^����x�w�].���v#����d)�u�}����w;��s9��W�U�u:=/�B ���L#���I$2����c�X��S�T
%���Z�F�`����f����`�t�m���~�G��h*5-��j��E�q�|����}�?���s9.�[-��j
���d��J�P�r�L����J�B����@  08<>��o���v�M&3�f	"�X&�Y,6;��s�\��s9.7�M�s��N�C�P��R����`(4��~���s�\�g�Y,�{=�o7���a0�����s9����u:=��k5��K%�i����W+
�����I����V��A 08<>������~�@����D��H�b�H�b�H"1,6�]����~�O'�D!�t�m��}��?�O�S��J�����H�b��D�a0�|��w;'�������I�r�s9�n����h*5-+�J���D�����A 0�|�o7�M�s9�w�].���v�M&�Y��[�������V�E"�X��S)���]��{=�o7�Q(4�}�����w;�N�C!�h�u��~����y<>?��g3��S)�u�����w;�g������r&3�L#��D��H"�X�f�I$���^�����@����D�a�x.���v����i4��~��g��l+�e2���G��h���]��{=�o���v�Q(��]�w;�g�Y��[��K%����M�s9�n�K��I�r�f	�b���B�`(��].7���S)�u:=��k5���[�V����P$��|��w;�N����@  ��\�g���V�E�q�|�o7��C�P��R��B��P��R	"�X&���V�a0�|�������W+
%�i�����k�Z#���l�k���f	"�X�s�\��s�\���t-+�J���`�t�m���~����D����L�c1�l�U*5������l+
%��J!����E�q���O��i4:=��k��M��y<>?�O'�D�a0��^�G#�H"�X�f	"�X&3��F��`(4�}����w;���c�X���i4��~�����|/���������`�h*5�m6�].��m��}��_/�E"�X�s9���}��_/�E"1���K%)��U*�Z�c�X&3���i�z�N��@  0��^��c1�l�k5�V��A�p�l��u���_/�B�@�`�h���]�w�].�[�V�E"1�v����p�v��C!(��].�[-����].7�M&3��y<>���w�]�w���W�U����n�K�R�D�a0�|�o7�M&3���|/�E��x.7���S)��z���c���F�A �x�����z��i4:�������^�G#�H"��L��h��U*5�m�{��O��i�z�N �p�v��f��d�i4�}>?����y<>��o�[-+�J��A�p��[�V�B��@�`�h*�Z��C�����A��X�f�I�����K%)��U��z'�D!�h*�����i���n�E��x��{���g3�L��q���O����Z�Q��Z��C�P���l+�e2�\����Z���a����G�Q��Z������L�Q(4�}�?�C��H��x���k5�m6;�N����H�b��D�P�d��J��p�v�M����^��a�����c�X�f�I���l�k5����m��}�?���@ �p,��}����������{=�o7���x.��m6������z��G���T��r&�����e29�n���r&����K%�T�e��|�o����[-�k5���e29���}>�_�W�U��z�����^���P��R	"���F���@����D��p�l�k5������[-��u:=��k���f�I�r�f�I�r��F������B  0�|�W��j��E�q8<>���w��n��p������������Y,������w�].�[-+��E���\�g3��F���P����d��t�m�����o�[��K�R���A�p,����_�W+���b�d)�j�J���D�����F��@��P���l+
����R	����T
%�i�z�N�@��P$�y�����{=/���r��F �p�l�k5�m�����o�[��K%)*��M&3����a�x�n�E"1��V��b�H��Q��Z�c�X�f	�b�H�b�H"�����a����G����J���`(�z�N�C!�t-��j�J�B��@  08�~�G#�H�b�H��x.�[-+
�R�D��p,6;�g3�f��d��J����P�r�f������R	�b��Y�����[�V����P��R	���h��U�u:=/����P�d���Z���x�n�E��x�n����Y,��}>�_/�K%���Z�F��@�`�h����U*5�m��}>�_/��A�p�l��u��~�O�S��J�B������@  0��^�G#�d���Z��C�P$29.��m6������z�N �p���K����R	�q8<���_�W�U�u�}�?���s��N�C��H�b����A 08��_��k5��v�M�s9��W+�e���^������F���H"1��[-�k5�m�{=�����~���q�|/��b$29���}>?�O��i4�}����w;�����x�n�E���\�g�Y�v��h*5�m��}>?�O�S)�j��r�f��B��@�`�h�j���Y,���~�C�P$�y���o��m6��n�E��x.���v�F�@ ��X����t���[-�����U�u�}>�_/��p��V�E�q���O�S)���]��{��O��i4�}>��������o7#�H�b����A 0��^����X�f��d�i�z�N���p,6;�g3�f�I$��|�W+
�R��B�@����D�a08�~�A�p�l+��E"1,�{=�W��j�e�y<>?��c1��V����P���I�r�f	"1��V���D�a08�~�C����B�`(4:��O'����`�t�m��}�?��c�X�f���R�D���X&���V��b$29�n�E"1�v�M&3�L�c�X����t�m�{=���u:=/���Q(�z��G#���B�@�����B�@�`�h�u:������|�W�U���]��{�^�C!��Z�F�A 0�����s�\'	���h���]�w;�g�Y,�{=�o���v#����A��X�f����I$�y<�������o��m6�������]���}>�_�W�U��z��s��N��`��T�e2�\'	���h��U*5�m�����o7��C!����f�I$�y����w;�N���p,�{���g�Y����v�F��@�`�h��U*�Z�F�@ �p�v���x��W+��E"1,�{=�W+��E�q�|�o7�M�s����c��L��h��U*5�m����_/�K�R��B��P$�y��_�����]�����_�W�U����n�K%��t��v�F�A��X&3��F���P�d�i4��~�O'�I$2��N��@������A ���N�C��H��Q�t�V��b����d��J�a0���O'������H�q�|/���r&3&3��S)����U*5���[-+�e�y<���o�[-����].��m���~��g��l�k��M&3���C��H"��L�c1�v�����X&�Y�v�F  08�~�O��i�z�N��a0��^��c�X�s�\���y<������w�]��{=�W+�J�B�`�h��z�N�@�`���J��p,�{=�o���v#�r�L���T
%�i�z�N��`�h*�Z�F  ��\'�D!(�z��G��h�j����Q��Z�c1,�{���g��l��u��~�C�P���I����V�B ��X��y<>��o�[-��u:��O'�D!����E"������p,�{=/���r����^�A����F�@  �������x��W�U*5-�U��z'	�b�d�i4:�^ �p,���~��g�Y,6��n�K%�i4�}���_/�P������I$��|�o7#���I$2���G#���I��Y,6;'	�q8�~�C��H�q���O��i4�}�����?��g3�L��q8�~�O��i��]�w��n�K���d��J��H�������q8<>?���P�d�T�e��|��w��n����h�j��r���C����B��������@  08<���?��g�Y���m6;'��d�i4:�^�C��H�b$29�n�B�@  0���O�S�T
�R������H��Q(��].���v��C!�t���e��|/��e�y�~��g3�L�Q��Z�c��L#�H���h�j���Y,�{=����z��G#����V!��Z#�H�b$������s9��W+�e�y<��?���q�|/����P$�y����w;�g3�L#�H"1��V!����E"���F���P�d)�����������j��E�q8<��_��������k5����m6��n��A�p���K%��t������[-+�J��p��[-+�e�y<>�_/�E"�X���i�z�N�C��H�q��^��`�t-�U*���f��B�@�`���J!����E�q������y<��?����y<>����{��O'��d�T���Y,6;�g���V�E���\�g�Y��[�V��A�p����v�����t�m6;�����x.7�M�s9���k�Z��h��z�S)���j���Y��[�������V�B���@  �x.�[�V��p�����r���C�P$29�w�].7�M�s9�n��b�H�q8<��_/�B��@ �p��V���D�P�d)���j��E"���F�A�p,�{=/��b����V!�h��U��z����q8<>?��g3������X�f�I$�y<>?�������O�S�T�e29�w�].���v�M&3�L�Q(4:=�W�U�u�}>�_�W+���Y,6;'�I$29�n�a0�|��w;��G�Q(4��~����y�~��a0�|/�K�R	��Q(��].7��f��B�`��T����l�U*5-�k5��v�F�A �x�n�K%�����f��B��@�`�h���].7��q8��_/����h*5-�k�Z�Q�t-�k�Z��C�P������������e��|/��b��D�a0���O'�I�r��S)��U�u�����w��n��e2�����q8<>���w��n�K����R������H"1,6�].���������v������Z#�d��t�m6;���c�X�f��d)*�Z#�H�b�H�q�|�W+�J�B�@���������H��Q�t�m��}>��o7��f�D�a08�~�G����J�B���@����D�P�r��F���H����������N �������p�l��j
%��t��v�Q���M&3&�Y,6�].�[-�U����n��e�y�~��g3&3�f�I�r�L#��R�D!���J���`�h*�Z��C!�����b���B�@ �p,�{=���{��O'��d��������t-��u:�^�G�Q����f��d��J�P$���^�G#�H"1�������l���z�N���@��P�d��t���[-����]�w;�N �p����v��q8�~��g3�f�I�r�f�D�a0��^�A�p��V��A �x��W�U�u����o�[-��j��E"1��V���Q(�z��G#�H"1���m�{=/���`����f	"��L�c�X��S��J���D���D�P�r�f�I��Y���m6�]�w�].7���a08�~�O��i����W+�J��A�p���K��I�r�L#$�y��_/���`�����b�H�������b����A�p,6;��G�Q(4:����s9��W+�e��|/���Q(��]�����_�W��j
�R��B�`��T��r��F�@  08<���?���p,���~�O�S�T
��I$29.7��h�u:=�W+�e��|�������o�[�V!�h��U*5�m�{��O�S)��U*���f�I�����K�R����`�t�V�E"1�v��f������H�b��D��H����N��a08<���o������v��q�|�o7����i�z�g��l����j�e2�\��i4���_���u:=�o7�M&3�L��q8��_/!��Z�F���P$�y�~�����|/��e2�\�g3������M&��l+
�R�������D��H��x.7����\�S�T
��I$�y<>��o�[-��u�}����_�W������j�e29�n�B����@ ��X��y��_�W���U*5�m�{�^�A�����C�P�d�i4�}>�������_���u���_/��e29�n�������K��I��Y,6�����u:��O�����M&3�����Z��h�j
%�T��r��S)���j�J����P�r���|�o7������b��D�a�x.7�M&3�f�D������������C��H�b��R	�����J�����H�q���O�S�T
%��t�m�{=�������o7���a�x�n��e29.��m6�]��{=������_���u:=/���Q���M&3��S��J�B�`(4�}�?�O'������R	��Q(4��~�O�S�T���Y,���~�O�S)�j�J���`�t�m��}�����{=�o7��C��H"��L���x.7���a08<��_�W+�e�y������}>�_/��e����O�S���E"����������C!(�z�N�C!(4������{�^����D�P��R�D��p,�{=/�E���\����|����}>?���q8<�?��g3�f��d�i�z�������g�Y��[���e���^�G#��R	�b�H"1��V�E"1��[-+���b����A 08�~�O'�I�r�L�c1��V��A�������p�l��u:=/����P��R��B�`��Z�c1�l��u:�����y�~��g3��F ���L�Q�t-�k5-+��E"1��[-+�J�B  ��\��s�\'����`�h�j
%��t�V�E�q8��_�W�U��z��G�Q(�z��G�Q��Z��h*�Z�c1�l��������u:�^�G#�H"1,�{���g3����a08<>�_���u��~��`(4�}>?�O�S����b�H��x.��m��}��_/�E"1�l�����n!�t-�U�u:=/��b������I��Y,6;����q8<>?�O'��d�����Q(���n��e�y��_��k��M&3�L�c�X�f�I$�y<>?����y�~���s9.��m6�]�w�]�w;'	"1���K�����I��Y,�{�^�A �x�����_��k5-��u�}>�_�W+�e�y<>�_/�B�`(4���_�W+������K���d��t�����v#���B �p���m6;'�I$2�\�g3&�Y�����[�V�E"1����v���a0��^�����L#�H��Q(�z��G#$2�\'	��x��W�U���]��{=/���Q�t-�����n�E�q�|�o7��C���D!(�z�N�@ �p����e���^�@  ���N��a��\��i4����o��m�{��O������f�D!��T��r&3�f	��Q�t-���z�N �p�l�U�u:��O'��B�`(�z�N�����B�`(4:��O�S)���������j�J�B�`���J��p�l��u:�^��c1��V�E"��L���T������K�R	��Q���M�s��N��@  �x��{�������^��c���F�@�`�h*��M�����O�S�T
����R	���h�j
��I$����O'���R	�q8�~�����D��H���h�u���_/�K�R�����P$2��N��`(4�}�����{=�o�[-+�J�B��@����D!�h�u�}>���w���������W��j��E�q�|�W��j
%�i4:���g3��F���@  �x������o�[�V����������P��R	"1�v�������M�s9��W�U*5-+������T
%�i4��~ �p,��}>��o7�Q�����S)���j�e�y<>�_��k���f�I$���^����x�n�K%��J��A�������p,6;��s��N�@�`��T
��I��Y�v�M�s����c1�v�����X&3�s�\�S)�j
%��J��A�p����v#��D��p,6�]���}>?�O'�I$2�\�S)�u:����s�\'�I$29.�[�V������D��p�v�c���F�A��X�f	��x�n����Y������m�{=��k5�V�E���\��s9��{�^�G#�r�L�Q(4:=�W�U*5��v��f	�q8<>?��g��l�U*5���e29�n�P�r��F���@�`�t�m�������{=/���Q(4�}�?�G�Q(4:=�W�U���]��{=/���`�t����m6�����u��~�G�Q(4��~�G����J�a08���o7�F��`��T
���d�i4:=/��e29��W�U*��M�s�����q8<>���w;�N��a08��_/�K�R	���h�u:=/!��T
%�������T���Y�v�F ��X�f	"��L#$2�\�S��J�P���I���l��u�}��?���s9���k�Z�c1�l�k�Z�F�`�t���[-��j�e�y�~��g��l�U�u�}>?��g3��S��J�a08<>?�A 08�~�O'�I$2�\�S��J�B�@��������P�r�L�c1�������l+��E�q�|�o�[-�k5��v�M��y���o�[�V�E�q�|���u��~�O�������������S)�j���Y,��}���?���s�\�����^�C!���J�a08�~�O�S)��U*�Z�F��`��T��r��S����b�H�b$��|�W��j
�R��B  08<>?�O�S)����U�u��~��@�`(4:=/����h�j
��I$29.7���x.7�F�A�p,�{���g����K%��J��p,���~��g3�L���x��W+
��I$���^��c��L��q8<��?  08<>?�G�Q�t��v�M�s9����~�C!(4����o7�Q��Z��q8�~�O'��B�`�h�j��r�f�D!(4:=�W+��E"��L�c1�����r�L�Q����f�����P��R��B ����F�@  ��\�S)�j
%)*5�m���~�`(��].�����m��}>?����x���k��M�s���G#�d�T
%�T
�R�D����L#���I$29�n�a��\��i4�}��_/��e2���G#$29.���v�M&�Y��[���e29.7�F���P����d�i��].7�Q(4�}>���w�]�w;�N�`�h��������z�����^��c�X���|��k�Z��C!�t-����].���v�F��P�d)*�Z����\�S�T����l�k5�m6��n��A 08<>?����D��p�v�����t�m�{���g3�f�D��p,6;���c�X&3�L����\'	�b���I$�y��_�W+
�R	"1���K%���Z�F�����D��p��V���Q(��].�[-�����n�������K%�i��]�����_��k5������[�V�P���I�r�L�c�����a0��^��c�X�s��N�A ��\��i4��~��g���V��p����e������s9��W�U*��M�����O���t�V��p��[�V��A 08����w�].�[-�k5-��u�}>?�O�S)�u:��O'�I�r�f	�q8<>��o7�M&�Y�v�Q��Z#$�y���o�[��K%����b��D�a�x��{=�o7����i�z'���R	�q�|�o��m�{=��k�Z����p�l��j�J�B��@��P���I�r&�Y,6��n���r�L��h��z����|�o7���S)*�Z��C��H��x.7����i��].7��h*�Z�c1����e���^��c��L�Q�t���[���e2����c1���K���d)�j���b�H����N�`��T
%)�u:=��k5�V�E"1��V�E"�X&3�L����\���t�V����h*5���[-+�J�B�`(4:�^��������a08�~�O��i4:�^����x��W+���b��D�a��\�g�Y���m��}>�_�W��j�e�y�~���p���K�R	����T
%)�����j�J��A 0���O��i���n�E"�X����^�C!�h�u��~�O'�I$�y<������o7���a0��^�@���H��Q�t����r�f�I$2�\�g3��F�A �x�n���r�f�I�r�L#�������r&�Y,6�].���v���a08<>�_�W+��E��x�n���r�L#����d����M&3��F�A 08<�?�A�p,6�]��{=��k5��K%)�u:=�o7�M���|��k��M����^�G�Q(��].7��C!(��].7�Q�t�m�{=�W�U*5�V!�h*��M������g3&3�s9�n�K%)*��M&��������l���U*�Z#�H�b�r�L�Q(�������z��G#�H�b�H��Q�t��K�������R��B�@  08��_��k5-�U*��M��y<>?���p�l��j�J��A�����C!�h�j�J!(4���_�W�����U*�Z��q8�~��g3�L#�d�i�z���c��������L���x�n���r��F ����F���H�b��Y�v�M&3���C��H��Q��Z��C!���J!������i��]��{=��w;��G�Q(4:���g�Y�v�M&3��F��`(4�}�?�O��i�z��s��N����@  ���N  ��\��s�\�S)�j�J��p,�{=��w�].���v��C���D!��T��r�L����\�g������r�f���R�D�a��\�g3�L�c�X�f�D!�h������U�u�}�?����x�w;��s9.�[-�U�u�}���?�G���T
%�T
%�i�z��G#$29�n��b�H��Q�t��v�c��L#�H��Q���M&3��y<�?�@�`�t�m6;����|���{=��k5�m�{=��w;'��d�T
�R	�b$�y<����w��n���r�f���A�p���K��I$�y<�����o�[-�U�u:=/��������e2����c�X�f��d�i4�}��_/��e2�\������������f��B�@��P$�y<>?�O�S�T
%�����f�D��p����v�c1�l��u��~���p,6;�����x�w;�N��a����G����J��A�p��V��A��X�f�D�P��Y,6�].7�M&3�L�c1�l��j
%)����n���Q�t-+�J�B�@ �����C��H��x.7��C�P�d)��U��z'	����N��a08<��_/�E�q�|�W+�J�P�d�T����l�k�Z��C!�t��v�M&�Y,��}>?��g�Y��[�V�E"�X&��l�k�Z�F���P��R	�q������y�~��a0�����s9��{��O��i4�}>?�G#�H"�X�s9.���v��C��H�q8��_/��e��|�o7�F�`���J�B���@�`(4:��O'���R	����T�e��|���{=�W����j����Q�t��K%)��U*5�����v�c��L��h�j�J!�h*5-+��r���|���{�^�G#�H��Q(4:=/�K%���Z���a08<��?�O'	���\�g3�f	"��L�c����C!������Q(4:��O�S)�u�}>?��g3����^���q��^�G#�����`(���n�E�q8�~�C�P���I$���^�C!�t���[-+��E"�X��S��J�a0�|/����P���I$�y<��_�W+�e29�n�K%)��U*�Z��C�P$2�����q�|���u������{=�o7�c�X������M���|�W���U���].�[��K%)�j�J��A �x��W+�e29��{=�W�U*5-�U*5-+
��I�r��������S��J����P�d)*���f�D�P$29.7�Q(�z�N�@ �p��V!����E"��L�Q(����W+�J���`���J�B�@ ���L��q8<>?�O�S)*�����i4���_�W+��E����N��a0��^�@  08���o7#$29���k5�V!��Z�F�A ����G�Q(��].���v�M��y�~�O�S��J����P�r&3&3��F��@�`�����b��D�P�r�f�I$���^�@  0�|/����h�u:=/�a���N��a0�|�o7���a�x�n�E"�����a����������G��h*��M�s9.��m6��n�E�q��^�G#�d��t��v�M����^�G#����A�p,6�].7�M��y��_/���r&�Y,6��n��e2��N�C!(���n��e2��N�@�`���J��A�p�l�U*������t��v���T�e2������x���k5�V�E���\'���R	"1���K%)�j�J��p�l�����n��H�q8<��_/����Y,��}������_�W+
%�i4�}>?�O'��d��J!������Q(�z��i4�}>��o���v�M�s9.7#�d���Z#��D�P$29���k5�m������w��n�K�R	��x�����z���t��v�F�A 08<��_/���r�L#��D�a0�|�o7�F���P�d��t��v������Z�F���P$�y<���?�C!�������t��v#��R�D!����E���\�������S���E��x.7���S)��z�����M&�Y,�{�^��`(4��~��g�Y��[���e2������x�w��n���Q�t-�����n�B����@����D!��T��r�f�D��p�����r�L����J!�h*�Z���x��W��j�J��A ���N�A�p,��}��?��g3�L#�d�����f	�b��D�a�x��W�U�u�}>��o���v�M&3��S�T
%��t�m��}��_�W+
�R�D!�t���e2�\��s9.�[��K�R	��Q(��].7#$���^�G#�����`���J��A 0��^�A��X�f�I�r�s9���k5-�k��M&�Y,6;�����M�s9�n���Q(4�}���_�W�U*���f�I�r���i4�}>�_�W+�J��A 0�|/�E"�X�f	���\'���R����`��Z��q8�~�����|���{=�o�[�V�B�@�������`�����b$�y��_/�K%������S��J!�h*5-+
��I�r���C�P�d�T
�R	�b$29.7#�r�s9.�[������l������W�U���]�w���W+���b�r�f	�b��D�a�x�n�E"1�l+��r��S���E�q8��_�W�����U��z'��d�T
%�T
�R��B�@ �����C��H�q8<>�_�W+���b��D���D�P$29�n�B��@����D!��Z�F�A����F��`�h*5-�k5-+����Q����f	���h*5�m6�]����~�G#�H���\���y<>��o7��q�|/�K�R	�b$2��N����X��y<>�_/�B�@�`��T���Y,��}>�_/�E�q8<��?�C��H��x�n���r���|��k�Z��q�|�W��j
%�i�z�N  �x�n������V!��Z�c1,�{�^�A �x��W���U��z�g�����e�y<>?��g3��F�����D��p�������l+���b�H���\�g��l�k�������Z��C���D�P�d�T
��I����V�B��@���H��Q(��].�[�V�E����N���P���l����j�J!��T
%)�j
�����I��Y,��}�?�G�Q��Z#����V��A �x.7�������Q(4����o��m6�].�[��K���d�������i�z�g3���C!���J�B��@���H��Q(4��~����y<����o7#�����R	�����J�B�@  �x��W+����l���U*�Z�F��@ ��X����^�����\���y<>��o�[�V!(��].������v�Q(�z���c1���m���~�G����J��A�����C!(�z��������G#��R���A��X��S)�j
%�i�z'���A������a�x�w��n�K%�T��r&�Y,6;'�I���l+��E"���F���P�����R	�b���l����j�����V�E"�X��y<����w�]��{�^�G�Q(��].�[�����Y,6;�g��l��u�}��_/���X�f�����d���E"1,6������z����q��^�G�Q��Z�Q(���n�K%���Z�c���F�@ ��X��y<>?�C!�h�j�J�P$�������y<���o���������v��h�u�}>?�G�Q��Z��C!��T
�R	�q�|��w�]�w���W���U*���f	��x��W�U���]��{=�����~�G�Q�t�m���~��g3�f���R���A��X&3���C!�h*��M��y<>�_/�K�R���A��X�����Z�F�@��P�r�s��N��a��\�g3��y�����{=/�P�d�T�����V���`�t-�k��M�s9��{��O�S�T��r��F���@ ��X&3�������L������G#���I$�y<>?���q�|�o��m6;��s9��W+��r�f	���h*5�V���X�s��N��a�x�n�B�@  08<��_��k�Z#�H����T���Y��[��K%)*�Z��q8�~�G�Q(4:�^�@ �p���K%��t�m�{=�o�[-��u:�^��@ �p��[�V��b���B��@�`(4��~�O'��d�i�����k��M&��l+�J����P�d����M&�Y,�{=��w�]���}�������_�W+������T
%)�u:�^�C��H"1��V���Q�t��������v�����t�m��}�?��a�x.����[�V��b��D�����F��P��Y,���~�O��i�z��s9.7����i4:�^�G�����E"����C!���J�P��Y��[�����Y��[-+
���d)�������u:��O'�I�r�s�\�g3�L���x���k5��v����p�l�U�u�}>��o7�M��y<>�_/�K%��������t�m6;������\�S)��������z�����^��c1��[�V�B�@�`�t�m��}�����o����[-��u��~�C!�t�m�{�^��c1��V!��T
%��t�m6;��i4:=�W+�����h�u�}�?���s9�n�B��P�d�i4�}�����w�]��{=�o�[���e29�w;��s��N�@�`�h���j�J��p��V!�t�m�{=��k5�m�{=�o7#�d��J�B  08<��?�G#�r�L�Q(4:=/�K�R�D!�t��K�R	�b��D��H��Q����f�I���l�k�Z�Q(���n�K������d)��U�u:�^�����L�c�����a0�|�o�[�V�E"1�l���z�S)�����j�J�a08�~���s9.7��f���R�D��H��Q�t�m�{=��k���f��d��t��v���S)�j�J�a�x�w���W+��E"��L�c��L#�d��t��v�M&�Y,����_/���`�t�����v#��R	��Q��Z���x�w�].7�����t�m�{������|�����~��g3���i4:=�o��m�{=/����L�����E"����C!�t�m6��n�a08<�����o7��f��d)*�Z�F�A ���N�A������a08�~�O'	����N  �x�n���r��F �p��[�V���Q���M&3�L�c1����e2�\'�I$�y<������o7�Q�t��v�M&3��S)*5��K%)*��M����^�G#�H�q8����w���W�U*5�m6;��G#�d�i�z�N  0�|��k5-��u�}>?�@����D�a��\��s9�����z��s9.7��f�D!����E"�X����t-�k�����i4:=/��e2��N�A 08����w;�S�T
�R��B�`��T�e29�n���X�����Z��h����U*5-�k���f����I$�y<�?�O�S)��U*��M�s9�w;�S������h��������U*��M�s�\������O���t�����v���a�x.���v��h���]�w;�g3���|����z�N�C��H����T
%�����f	"�X&��l���z�N�A��X�f��B�@ �p,6���W��j�e��|�o7��C��H��Q��Z��������C��H���\�g�Y�v���x��W�U��z���c�X&3�L#���I$2�\'��d�i4:�^��a0�|/�E�q8<���o7�M��y<�?�O'�D�a08���o�[-+�J�a����G#$29.�[��K��I���l�k�Z�F��@�`��Z��q8<���o7�Q(4:=�W��j��������r��S)����U*��M&3&�Y,�{=�����~�O���t-+
%�i��].���v���a08<���o7�F�A 08������}���_/���r���|��w;���t��v�c�X�f��d������S��J�B�@�`�t-���U���].7��f�I$�y�~�O'	�b��Y��[-+�J�B�@�`��Z�c�X&�Y��[�V�E"1��[-�k5-��j
��I���l��u����o7�M�s9���}>��o����[��K��I$�y<>���w;�g3����a�x��{=�o7����p�v�M&3&3�L��q8����w�].��m���~�O��i4:=�o��m���~�C�P��Y,6�].7�M����^��c1�l�U*���f��B  08��_/����Y,���~��c�X�����Z��h�j�e��|/�K�����I$2�\�g3��F�`(4�}>��o7�c1,6����k��M�s9���}��?�������O'�D�a�x.�����m6;'	��������Q(�����k5��v�����t��v�����t���[���e�y��_�W+�J�B�@��P�r���C��H�b�H"1��V���������Q���M&��l�k����S)����n�E"1����e29.��m6��n�K%�i��].7�c1�v�Q(4�}���_�W+�e��|�����~��c�X�f������H���\�g����K%����b�����`�h*5�m6�].��m��}>�_/�B  08<>�_/�E"1�l+
%�i�z�g���V�����H"��L���T�e2��N�A�p�l�k��M�����O'�I������e�y�~�����\�S)*5���e29�w;'�D!�h�j�J!�h���j�e�y<>?��a0�|/���`(�z����q8��_���u:=/����Y,�{������|�o7�M&3�f	�b�H��Q�t���e��|�W+�e2�\'�I�r��F��`��T
��I�r��F����H"����C!��Z��C!�h��U�u������{���g3�������L#�r�s9.�[��K�R��B�@�`�t���[-���U�u�}���_/�K%����b�H�����G��h�u���_/�����T�e�y<�?����@�`�t-+�J���X��y���o��m��}��?������N�C�P��������R��B��P��Y�v���S)��z�������S)�j
��I�r�L#�d���Z#�H"������p�l�������U���������]�w;'��d)����U�u:=�o�[-+�e29������].7��C!�t��v�c1�l�k�Z�c��L#��R���A����F������A��X&��l���U*���f	����T
��I$29.�����m��}>�_/�K��I$29.7�c�X��y�~�G��h�j�J�P$��|����}>?������N����@  0��^�A�p��V�����F��@  08<����_��k�Z�c����C!�t-���U���]�w�].7���x��{=�o�[-�U*�Z��C!���J�B���@  �x.7��C!�h���j�J!�h�j���b�r��y��_���u����o�[�V�����T�e�y�~����y����w�]�w�]����~�C��H�q8<>?�O'	�b�H"1���K��I���l+
%�i4:=�o7���a0�|�W���U*�Z�F���P$29��{��O�S��J��p���m6��n�a0��^��`��Z�F�A 08<>�_��k�Z��h��z'�D��p��[��K%�T
%)�j
�R	��x��W+��r�L�c1����e�y�~�A 08���o�[�V�E��x�w�].7��f�I$��|��w�].7�M��y<�?����x������].7�M��y�~�O'���R�D!(�z��i�z���c1��V�E�q8<>�_/�E�q�|�W+����l�������k�������Z�Q(��].7�c1���K��I�r�s9�n�E"1��[-+�J��A�p,6�]��{��O����Z���a08���o7����i4�}>�_/���Q(����W����j��E�q����g��l���U*�����i4:�^����X�s9�w�]��{�^�G#��R	�b��Y,6;����Z��C!�t�m��}�������_/��e��|/���r���|�W�U*���f��B  ��\'����I�r�L#�H�b�d���Z#$29.7�M���|/�K%)*5����r�L���x.�[�V��b$2���G�Q(4:=�W+���b�H���h�j�J��p��V��b�r�s9.7�M&3���C����B�`�h*�Z#�H��Q�t�V!��T
���d�i4����o7�F��`��T��r��S�T
%������h�j��r��S)���j�e29�n�K�R	�q����g�Y����v�M&3����a�x.7��f�I$�y<�?��g�Y���m6;�����x.7����p����e29��W�U��z�N�C!(�z'��d�i��]�w��n�K%)�j�J���`�h��z��i����W�U��z����q8<>��o�����m6;�N�@����D!���J���`(����W�U�u�}��_/�K%���E���\�g�Y,��}>?�O'�D�a0�������|/��b�d��t����m��}>?��c1�v��f	�q8<>�_/��b�d��t��v��f�D��H"1�l��u:�^�G�Q��Z�F�A��X����t�m��}>���w;�S)�u:�^���p���m6����k5�V���Q(���n���Q(�z'	"�X��y<>��o7���S�T
��I$�y�~��g�Y�v�M&��l����j�J�B  0�|/�K����R�D�a��\�g3�L#����A 08���o7�M&3�L���������x�n���r�L#�d�i�z'�I$2�\��s�\�g3�L#�H���h*�Z�����X���|/�K%)���j��E"�X�f	"�X���|��w�].��m���~�G����J���`(�z����|�o7��f	�q8�~��g����K�R	�q����g�Y,�������{�����y<>�_/�E"�X���|��k�Z#�d����M���|/��e29��W��j
�R���A��X�f�I$�y<>��o�[�V���X��S)�u���_��k5�m6;�N����D��p��V�a�x�w;��i4:�^�����\�g�Y,�{���g3�L�Q(���n��e29���k5�m��}>?�G����J�B���@��P��R�D!�h��z�N�A�p��V��b�d)*5�m����_��k5��v�M&�Y,6;��G#�H���\��s�\�S�����Q�t����m6�]�w;���c���F�@��P��Y,6;�N�A ���N��a08<����o7��C!��T
��I�r��F�A�p���K��I$29���k5-���z�N�@����D�a08�~������@  0����g3��F��`�h�u�}>���w;���c1�l�����n�K%�i4:=/�E"���F�A 08�~�O'�I�r�L#���l+�e29�w��n�K%��t���[-�k����S�T
%����M��y<>���w�].�[����r�L#�H���h��U�����W+
������d)����n�K�R	�q8�~��g3�f�I�r�f�I�r��F�A�p�l�k5��v��f��B�@ �p,���~���s�\���y<��_/�E�q���O�S)��z���y<�?��a0�����s9.���v�M&������r��y��_/�K%�T
�R	��x�w;�N�@��P��R�D��p�v�M&3�L#$29�n�B �p�v�F�@��P�d�i4:=�o�[�V�E��x.�[��K%�T�e�y��_�W�U*��M&��l����].7��f	�b����d�T
%��J����P�r�L�c�X�s9�����z�N�C!���M&�Y����v#���B��P���l�k��M�s�\�S����b�d�T
�R	��x������]�w�].7�M&3�L�c�X������M����^��c1�v��f��d�T
�R�����P��R	�����G#��D������`�h���j�e2�\��i�z���c1��[�V����h�j�����h�j�J��A�p��V�E�q�|��w��n�E"����C���D�P$2�\���y<��_/�B�@  08<>���w������z�g��l�k�Z�F�A �x�n���r����a����G��h���j�J�a0�����s�\��i�z��G�Q(4��~�G#�H�b��Y����v��C��H�b�r�L�Q(����W�U*������t�m6��n��e29�w��n�E"��L�c�X�s����c��L����J����L#����A ��\��s�\���t��v�F����H"1,6���W+
%��t�V�B�@ �p,6��n�K%��J��A��X��S�T�e�y�~�����\�S�T
%��t��v�M���|����}�?�O�S�T�e2�\�S)*5-�k5�m6�].�[��K%��J���`(4��~��c1��V����h���j
%)*���f�D!����f�I$�y<>?����y�~�G��h*5��v��C�P������I�r��S��J�a08���o7����p�l�k���f�I���l�����U����n�K%�i��].7�c1��V�E���\�g3���|/�K%)�j���b�H�b�d��t�m�{=��k5-+���b�d�i��].7��f	��Q���M&�Y��[�V�E"������p�l�k�Z�F��`(4�}���_�W+�e��|��w�].���v��f��d)�j�����V�B������A 08<>��o7���S)*�Z#������e�y�~�O�S����b�d)�u�}�?����y<�?����y��_���u:=�W�U�u��~�G��h�u:=���u�}��?�O�S)�u�}�?�O'��d�i���n��H��x���k5��v��f�����d���Z#�d�i4�}>?����y�~�O'	�b���B�����B��@�`���M�s��N�C!�t�m�{=�W�U�u���_/����Y,6;�N���@��P���I���l����].��m6;'��d)�u:=��w;���c�X��S��J�P$�y�����{=�o�[-�k5����r����a08��_�W�U*��M&3�L�Q��Z�c1�����r�L���T
%�i�z��s��N���p������m��}>�_�W+��E�q8<����w�].7��f�D�a��\��s9.��m6�].���v����i����W+�e������s�\���t����m6��n�K���d�i��]�w����k�Z�������c���F���P�d��t���[�V���X�f�I$2���G#�H"1��[��K�R	���h*5-���z�N�@�`�h*5�m��}����_/�E�q8<�?�O'��d�������i��].7��f	����T
%����M&�Y,�{=��w��n��A 08�~�O'�D�P�d�T���Y�v�F  ���N�C!(4:�^�G#�H�q�|���{�����y<���_/��b�H�q8<>�_/���Q(4:�^�G���T�e�y��_�W�U*�Z#�r�L#��D����L�c1�l+
%�i���n�E�q8<>?�C�P$29�n�����F�@�`�h�j��r�L��q����g3��F��@�����B  �x�n�K���d�T
%�i����W+
%�T�e���^��`��T
�R	�q8���o7��f	�b�d)�u:=�W+�e�y��_/�K��I�r�s9.�[-��j
%)�j�J�B���@  ��\�g�Y,6���W���U�u�}��_/�E�q��^�A ����G#�d)�u:�^���q8<>�_/�E�q8�~�O'���R	"�����a0�|�o�[-��j�J!����E��x.7��C�P$29��W�U*5��v��C!�h���j��r�L�c1���m6;�N�����L�c�X�f	��x�w;��G���T
%�T��r����t-+�J�����H���\�S�T
���d��t�m6;�g���V���X�s9.��m����_��k5�m���~�O�S)��U*��M&3��F�A�p���K���d)�j�e29���}>�_����z��s�\�g�Y,6��n�K�R���A�p�l+������T
%�i4�}���?�O'	�q8<��?�O��i4���_/�B���@�`�h��z��s9.������v�F��@��P$2�\����|�o7����i��].�[-+
%��J�����A 0��^ �p,�{=�W+��r����t-��u:=�o7�������M&3�f�I������e�y<��?��g3�L�c���F��`�h*����S)��U��z����q�|�o�[���e��|�W+����Q�t�m6�]�w;�N��a08�~�����|��w�].�[�V�B����@  �x��W+�J!�t�m���~�������O'��B��P�������d�i4:=�o7��f��d)�j�J�a0�|��w;�g3���C�P���I�r��S���E"1�v�M&���V���X�s9.�������[-�k�Z���x.7#$29�w;������\��s9.��m��}>?��g3����t��K%���E�q8<����_��k�Z�F����H��x��W+���b�H����T�e2�\�g��l���U*�Z��h����U����n�K%��t��v�F �p��V�E�q8��_�W�U�u�}����_/��b�H���h���j�����h*5�m�{��O'��d��t�m6�]�w�].���v�����X&���V���`�h�j��E�q8�~�O'	�b�H"�X&3��F��`��T
��I����V�B�@  ��\'�I�r�L�c��L�Q�t�V��b���B��P�d)��U�����W+�J�����A 0�|/�E��x��W�����U�u:����s9���k5-+�J�����H�q8�~�G#��D��p���K�R�D!�h�j����Q(4:=/��b�����R	���h��U���]��{=���{=��w;���t�V�B �p�l+�e��|�W+�J�B  08��_���u�}�����?��`���M&3&3&����K%�T
%�i4��~�C!(4:�^�������C!�t��v�M&3��F����H�b�d�T��r����a�x�w�]��{=�o7���a���N���p����e2�\��i�z'�D!�h�u:�^���p,���~�G�Q�t��v�M��y<����?�C!����f���R	"1,6;�N�C!�h�j���b��D��p,6;�S��J��A �x���}>��o7���T
��I$2�\��i4:=/!��T�����V����������������h�j�J���`�h�j�J�a08�~��`(4��~�O'�D����L�Q�t�m6;��s���G#����A�p,�{�^�G#�r�L����J��A�p�v#��R�D��p��[��K��I��Y,6�].7��q8�~��a08<>�_��������k5�m6�]�w��n�B ��X&3�����Z���T��r�f��d�i4�}��_�W+��E"1�l�����U*�Z����p�l�k�Z�F ��X�f	��Q����f�I��Y������m���~�O�S)����U�u:=��w�]�w�].���v�M�s9��W+�J�B�@��P$�y����w;���c1�l��u:=/�K�R	����T��������r����a08��_/�E"1�l���z�����^�`����E"1���K�R	"��L#���B�@  08<>�_/�K�R	���h*5������[�V�E"1�l������W����j���b��Y,6�].7��f	��Q(4��~���q���O�S��J�B�@�`����E�q8<>?��@  0��^�C����B�@�`�t���e���^�G#�r�s9�n������C!��T���Y,�{=��w���W+����Q(����W+�e��|/�K%)*���f��B�@����������D�a�x.�[-�k�Z�����N��a0�|��k5��v�c��L#�H"1�v��h����n�a08<>?��g3���i4�}�?�O�S)����U*���f��d)�u���_/�K%)�u:=�W+��E"1�l�����n�E"1��V����P���I�r��F�A ��\�S�����Q(4:=��w���W+�J����B�@�`��Z��h��z��G�Q(4:�^��c��L�c���F��@�`���J�B  ���N�C!�����S)�j�e��|��w���W���U������k��M�s�\��s9��{=�W+
��I$2���G#�H��x��W�U*�Z��C��H�b�r�L#$�y���o��m6;�N�C��H���h��U*5�V����P�d)�j����Q(4:=���{���g�Y,��}>?���p�l�k5�m6;�N�A�p,���~����y������}�?���s9�����z��G�������Q�t�m6��n��b$29��W+�J��p��V��A�p�l�k�Z��C��H"1�l���z�S)���j�J���X��S)��z���y<>�_����z��s�����q8<�?�O'�D�a08<������w�].7�F�A��X���|/�K%�i�z'	�b��D�a0�������|/���Q�����S�T
%)*5���[-�U*5����m�����o7�M�s��N�C!(4:=�o7����i�z'�D�P������I$�y�~���s9�w;'	��x�n��e29�n�������K%�i�z��G��h���j
%��t����r�L#��Y,����_/��b�d�i����W+
%��t��K%�����Q�t���[�V�E"���F�@  ��\���y<>�_/�K�R	"1,6;����Z����\�S)�j��E��x�w;���c���F��P���I�r���C!�h���]�w;�N�����L��q���O��i�z�N�C�P�d�T���Y,6�]��{=�W�U*5-��u:=/��e29�n����Y��[�V��b$2�\'����I��Y����v#��D�a08�~�O'��d��t�V��b�H�q8<���_/!(4���_/�E"����C�P$2�\'	���h��U*5-�k5-���z��G#��R�D��H"���F���P��Y��[-+��r�f	�b��Y,6;���c1�����r��S)��U�u��������~��g�Y,6��n�����T���Y,��}����o�[��K�R���A����F�@  0�����s�\'�I�r&��l�U*�Z�c1,���~��g�Y��[��K��I�������r�L���x���k5�m������w;'�D�P�r�f��B  08��_/�����l�U*����S�T
%�i���n���`����E"1��V�B���@��P��R	����T�e�y<��?���s�\�����^���q8<>������~�@�`�h�j�����h������U*5���[�V���Q��Z#�d����M�s�\'�I�r�L#��D�P$��|��w�].�[�V�E"1�l+
%��t���[��K��I$2�\�g��l�k�����i4���_/���r��S)���j�J!�h*�Z��C!�t�m�����o7�c1��[�V!�h*��M���|���{=/�����������l��j
%��J�a0�|�W����j�J������D��p��[-��j��E"��L#����A�p��V��A��X����t�V�a�x�n��e�y<���?�����L#���B  0�|�o7�Q(4�}>�_����z��s��N��@���H�b��R	����T
%�i4�}���o7�F�A��X�f��d����������b�H"1�l���z��i�z�N�@  �x�n��e���^�C��H���h�j�J�B���@ ��X�s���G#�H��Q(�z���c1,6;��s��N�C!(4:=�W�U�u:�^���p,�{=��w;�S�T
������d�i��]�����_�W+�J��p��[�V�E�q8��_/��A 0�|�o7�M�s9.����[�V�B�@ ��X&3&�Y��[-+��E"1��[-�k�Z�F����H���h�j��r��F���P�r�L���������x��{=���{�^�G�Q�t�m6��n���X&�Y����v��q�|/���r��S)�j
�R�����P�d�i4���_��k5�m�{�^�A�p�l��������u����o�[��K�R�D�a�x��W�U*5-�k�Z�F���H"1�l�U*5-�k�Z���a��\����|�W���U*��M&���V��A����F�����������@ �p,6�].7�M�s9�n��H�b$29�����z��G�Q(4���_�W�U�u:=�o7�Q(4�}��_/�K%����M��y<�����?��g3�f����I�r���|���u:�^�A 08<>�_�W+
%)�j
�R��B�@  ����G�Q(4���_/��e29��W+�e2�\�g3����a08<>�_����z�����x�w���W�������U*�Z��C�P�r&���V��p�l+�J!��T����l�k5�V��H��x���}�������_/�E"1�����r&�Y�����[-�k5�m6;��G#�d)��z�N�C��H�b�H"��L���x�n!�t��K�R���A ��\��s9�n�K�R���A 08�~�C!(4��~�O'	�b�d�i4�}>?�C�P$29�n��e�����g3��S��J!(4��~���q��^����x.7�M&3���|�W�U*5��K�R	�b��Y,�{��O'������H�q8�~�O'	����N�A���L����\��s9��W+��E�q8��_/�K��I���l��u:�^�G#$�y<>?����X��S)���j���Y��[�V���D!����E"�X&3&3���C!��T��r�f�I�r��F�`�h*5-��u:=����z��G���T
%�i�z���y<�?�G�Q(����W��j��E"1,����_/���r��y�����������{����s9������o���v���x.7�����X��S)�j��E"1�l�U��z����q�|�o�[-��u��~��������`�h��U*���f����`��������T
%��t-�U*�Z�c��L�c1��V�E"1�l����]�w��n�K%�i�z�N�C��H�q8���o�[-���z��s���G#�H"�X&3����t�����Y,�{=/�E�q8<��_/�K���d)��U*�������Z��q8�~���s�\�����^  �x��W��j
�R���A ��\��i�z��s9��W�U*�Z�F���@�`(4:���g�Y,6;'�I�r��y��_/��b��D�P�r�L�c�X&3��S)�j���b��D�P�d���Z�c�X�s��N����H�b�d���Z#���B�@��P�r��S)���j�e29�n��e2�\���t��v�M&��l�U���]��{=��w;�N��a�x.��m6;��G#�H�q��^��c1��[-��u�}��_/���r�f��d��J�a�x�n��e��|�W��j��E���\���y���o�[-���z��s��N����X�f�D�P�r��S)*���f	�q8<���_/�B�@��P��R	"�X&3���C!�h�j��E"�X�f	�b��D!�t��K�R�D��H"1,6���W�U*�Z#�H�q�|�W��j�J���`���M&��l��u���_�W+��E"�X�f�I��Y,6����k�Z�Q(4:=�o7�M&�Y,6�]�w��n��e29.���v����p�l��u:��O'��B��P�r�L�c���F����H������E�q�|�o7�M�s�\�g3�f�D!�����S���E"�X���|��w�].7��f�D�a��\���y<>�_/����������h*�Z���x��W+�J�a0���O'�I���l+�J��A�p�v�c1���K%�i4��~�O'	���\'��d�i�����k5��v#���B�@�`�h��z�N�A���L#�H�b�H"��L�c��L�Q(�z�N�C!�h�j����l��u��~�`��T
%)���].7��C!�h�u:=�o�[-�k5-�U�u:�^���q8�~��������a��\�S��J�B��P$�y<>�_�W+��E�q8<����o7����i�z��G��h��U*��M&3�L�c1�l�U*�����i�z���c�X��y<>��o��m�����o��m6;�S��J�B�@  ��\�g�Y��[-�U*�Z�F�@�`����f	�b$2�\��s���G#�r&��l����]��{=/�E"1��[-������j�J���`(�����k5�m6�]�w;�N���p���K��I��Y���m6���W�U*5�����Y,��}����o7�c1��[-�k�Z#��D�a0��^�A 08���o�������[-��u�}���?��c1����e���^�C��H����T�e29�n�E"�X��S����b$���^����X&3��y�~��g������r�L�Q�t��v��q�|/�K�R���A�p�l����].�[���e���^����x.��m6;�����x.7�c1��V��b������I$��|�o7��f��B����@�`�h*�Z�F�A �x�n�K�R����`��Z�����X&�Y,6;�������S�T
�R	"������p,��}���o�[�V!(���n���`�h����U*�Z�F��`(4�}>?��`(4:����s�\��s���G#��Y�v�F�A�p,6��n��b�H�b�d�i4�����w;��s9�w;'�����d�i���n�K�R	�q��^���q��^�����D!��T
�R	��x�w�]������o7�����N����H�q�|�o7�M&�Y,���~�G#��D���D!�h��z���y<>���w�].�����m�{=��k5��K�����I$29.�[��K�R���A��X��y<��?�O�����M&�Y,���~�C�P$�y���o7�F�@ �������p,�{=/���X&3��F�A 08<�?���s���G�Q(4���_/��e29��W+�J��p�l+�J�a��\���y<>�_���u��~�G����J����P��Y,6;�g3�L�c1�v�F��@ �p�l�k5���e29��W��j��r��F ���L����\'	��Q��Z�c�X�f�I�r�f��B��@�`(4�}�?��g���V��A 0���O'�I���l�k5��K��I��Y,��}��_�����]�w��n�B�@��P����V����h�u:=�W+�J����L��h��U*�Z�F�A 0�|��w���W�U*�Z����p��V����L�c1,6;�N��a08<��_�W����j
%��t��K%�i4:=����}��_��k5��K%��J��������A 0�|�o7���S)�j�e�y<���?��g���V!�h���j�����h�j
����R���A�p��V���Q(4�}�?�����\�g���V�B  �x�w;��G#��D��H���\���y�~�G�Q(4:�^��c�X�f�D!��T��r�s9�n�K%�i�z'�I��Y,6;���c1,�{=�o����[���e2��N���p��V�a�x����u:=���{=���u��~�G#�d��t��v�M&�Y,6;���t-�k5�m6��n�K%���E�����G#�r&3&3�L�c�X�f����I$��|������_/�E"�X��y<>���w;������\'	���h�j
���d)*5���[-��j���b�H��Q(�z��G#������e29.�[�V����h*�Z�F���P$29.7�c��L���x.������v�M&��l�k�Z���x�n!��T
�R��B�`��T
��I��Y��[�V��b��D��H���h*5�m�{�^�A����F�A 0�|��w;'�I$2�\�g3�L#�H�q8<>��o���v�M&3�f�I�r���������C!(�����k��M�s9�n�K�R	"�X�s9.7��f	�b�d��t�����Y�v���a0�|��k�Z#$�����g3�L�c1�l+�e�y<����o�[��K%��t��v����i�z��G�Q(4��~�O�S�T
���d�����f�I�������r&3&3�f��B�`(4�}�?��c1�l�U��z�g3���C!(4:�^�C!���M&3�L�c1�������v��f�D!(�z��G��h��U��z�����M���|��k5�m��}>?�O�S)�j�e2�����q8<>�_��k5�V������J�a0����g���V��b$2���G�Q���M&3��F�A 08<>?�O�S�T
�R��B�@�`(��]�w���W+��E"1,6��������n����P�r��F  0���O'��d��J��A�p,6;�g3�L�c1��V�E"1�v��h���j�J!�h��U*����S)��U*��M��y<>�_�W+�e29���k�Z�F��P���I$�y��_���u:���g3��S��J��A�p,6;���c1���K�R	��Q(��].�[�V�����T
%�T
��I$��|���u:����s9����u:=��w;��G�Q(4:�^�G��h*5-�������k��M&�Y,6�].����[-+�J�B�@ ��X�f�D��p��V�a��\�g��l��u�}>������~�G�Q(4:�^�G#���B  �x���}��?�G#$����O�S�T
�R��B  ���N���H���\���y<>?�O����Z#�r����a08<��_/�K%�i4:�^���q�|�o�[-�U*��M����^�G��h�u:=��w�].��m�{�^���P$2�\�g3&3�f�D�a0��^�����D���X�s�\��s9.�[��K%�T
%)�j�J���D���������X�f�I$�y<>?�G#��R	�b��D��p��V���Q�t�m6�].����[-�k5���[-+�e�y<��_�W+
�R��B�@  ��\'��B��@  0�|���u:=�o�[-�U*��M�s�\�S)*5�m�{��O�S)�u�}>�_/�����T���Y���m����_�W�U*5��v���S)����U�u�}����o7���a0���O'��d)*���f	�����J��A 08���o�[���e2���G���T
�R��B  ��\�g3�s��N�C!��Z���T
���d�i4��~�O�S�T����l+��E�����G#�H��Q(4���_/�K%)*�Z��C����B�@  08<>?��g��l+�J���X����^��c1���K%��t����m6�].7��C�P��Y��[�V������`����E"��L�c�X��y<>?���s9���k5-+
��I$2���G���T
%)��z'�I���l�k5-�k5���[��K�������R�D�P�d�i�z�N��`�h��z�S����������b��Y��[-�U*��M��y<>�_/���r&3�s9��{=�W+�J�a08���o���v����p��[-�k5��K��I$2�\�g3�L�c��L���x����~�O'�I�r�s9.�[-�U��z'��B����@ ���L�Q(�z��G#��D���X�����O�S)��z�g3�f	��x.�[-+
%�i��].7�����N�A 08<��������{�^��a��\��s9��W+
%��t���[����r&�Y�v����i4�}�����_/��e��|�W+
�R	��x��W+
�R���A��X��S)�j���b�r�L���x�n���r&�Y�v#�H�b�����R�D�a08<�?��������g��l�k5�m��}������}�?����X����^���p���m6�]�w;��G�Q(4:�^�G#��D!���J�B��P������I$2�\������f��d�i4�}�����{�^�G#�����`(�z��i���n�B  �x�w��n�B�@��P$��|����}>���w����k�Z��C���D!�t�m�{���g��l��j��E"1,6�]�����_�W+������������T��r&�Y,���~�O�S���E"1��������[���e2�\�g3�����p�v�M�s��N��`��T��r��F����@ �p,6;�N�C!����E"�X&�Y���m����_/�B��P$�y�~�G#�H��Q(4:��O���t-���U*���f�I�r���i���n����L��h���j�J���`�h�u����o�[-�U�u:=�o7�F�A���L#����d�i4�}���_�W+
�R	"�X���i4:��O���t�m�{=�o�[��K���d�i�z���c�������X&3�L�c1,��}>�_/�E"��L�c���F  ��\�S�T
�R	�q��^������N��`(�z�N��`��T�e����O��i�z�g�Y��[�V��b$2��N ����F�A��X�����Z�F  08<>����{�^���p�v��C����B�@ ����F��`(4:=/�����H�q��^��c1�l�U��z�N�@  08�������~����x���k5�m���~��g�Y,��}������_���u:��O'	�����J���X&3��y<>��o��m6;�N�A ��\'�I$29.�[-�����n�B�@ �p���K��I$29�n��A ��\�g�Y,6��n�E"��L�Q��Z��h��U�u��~�O'���R��B���@�����B ����F�@�`���M��y<>?�O�S�T�e2���������G��h*5�m�{�^�G�Q(���n��H�b�H�b��R�D�a�x��{=�o�[�V�B��P��Y�v���a�x���k5��v��h���]�w��n�B�@�`(�z�����x�n�K���d�i4:=��k������t-����]�w���W���U*5-��j���b$2�\�S�T���Y,�{�^��a�x��������{=/�K%�T������K�R�D!����f���A �x.�[���e�y�~�����L�Q����f�D��p�l��u:��O'��d�T
��I$�y<>?�O'��d�i4:=/��A�p,�����o���v��f���R�D�a0�|�����~�O��i�z�N ��X��y<���?�C!��Z�����N�C!�h*�Z��C���D��p,6�]��{=�o7������L�c1�l��u:=/�K%�T
����R����`����f�D��p�v�F����@ �p,�{=/������V��H"�X�f���R�D���X&3�f	�b��D���X&�Y,6���W+�J!(4:�������^�@�`(�z�g���V�a08��_/�a0�|������n�E���\�g�Y,��}>��o���v����p�l+�e�y<�����_��k5-����].�[��K%)���j�e�y��_����z'	�b�H�b�d)���]��{=/������V�B ��X�����Z�F�A������a����G#��D��p������Y,����_/��b��D���X&3��F�A�p,��}�?��g���V�E�q8<>?��`�����b�H��Q(4:=/�K%�i�z�N�A�p�v������Z�Q(��].�[��K�R	�b����V�E���\'	�b��R�D�����A��X���i���n�K��I$2��N�A 08<����o������v��f�I������e�y<�?���s��N�C!�t�m��}>�_���u:�^��`���J!(��].7���T��r&�Y���m6�].�[�V�E"�X�f��B���@  08���o7��q8�~���s9��W�U*5�m���~��c1�v#�d)���]�w;'�I�r�f�I$2�\��s�\��s����c�X��y<�����_/���Q����f�D�����A ��\�g�Y����v�F  ���N�@��P���I$��|�o��m����_�W�U*5�V�E�q8��_/�B��P$29.7�c1��[�V�a08<>�_�W�U���]��{����s�\'��B����@ ����F��`�h��U��z��G�Q�t�m6�]��{=��w�]�w�]������o7�M&��l��u:=�W������j�J�B�@��P���l+��E�����G#���I��Y,�{��O���t���[��K%)�u:�^��@  �x��W�U�u��~  08��_�W+�J��A���L��q8<������w;���y<>��o��m6���W�U*5��K��I���l�k5�����v��f���R��B��@�`�h��U*��M&�Y,6�].7#$2�\�g3&3�s�\�g3��F��P�r�L���T
%)��U*5�m6;'���A 08<>?��c��L��q8<>?�O'����`���J�a08<��?�O'�I$29�w���W��j�J�B����@�`(4��~��a�x�n�K�R	"1�l��u:���g3&3�����Z#�d)���j
�R	�b��D�a�x��W+�e29�n��H"1��V��p�l���z��G����J���`�h���j�J�P$29�n!(���n��������e29�w�]�w��n��e�y��_�W���U����n�K%�T
��I$�y��_/���Q(4:=/�E�q8<�?�C��H��Q(4:=/��e����O'�����d�T
�R	�b���B��@��P���I$29�n�B ���L#�H���h�j�J!�h��U��z�g3�L#$�y<>?�O��i�z�N��a���N�C��H��x.7�Q(4:=�o7�M&�Y�v�M&3�L�c1,���~���s�\'	�q8�~�G�Q(�z������\�g��l������j�����h�j��E�q8<����o��m6;�������g3�f�D���D���D��p�v����p,6;���c��L����\'��d�i�z��s9.7��q���O'�I�r&3��S)��U�u:�^�G#$��|������_��k��M���|�W+�J�B��@ �p�l�k5-�k�Z�F��`���J�a�������x�n�K%�i4:�^��c�X�s9.7���S�T�e��|�o��m6;���y<�����o�[�V��A 08<������_�W+��E�q�|�o7�F��P��R��B��P�d�i��]���}>?�@ �p�v�M���|/����h��U*���������f�I��Y,6;�S�T��r�L#����d)�j���b�H�q8<���o7��f������H"��L�Q(4:=�o7�c��L�c�X�f�I�r���C!�h��z��G#����d�i�z�����x����u�}���?����y<���?�O'�I$�y�~���q���O'	�b�d��t�m������w;����Z�c�X�s�\'�D!����E"1�v#���B ��X�f	"1,�{=�o7����i��].�[�V������D!��Z����J���`�h�u��~��c�X&���V��b�d)�j��E"�X��y�~���s9�n��A 0�����s9�n�K�R�D��p,��}������w��n�E"1�l�k5�V�E"�����a0��^�G�Q�t-���U*5�V��A 08<>�_/�K����R��B�`���M&3�L��h*����S)*5�m�{=�o�[��K��I$29�n��e��|��k�Z�c��L#��D!���J!�h�j
�R	��x.7���S)��z'���R	"1�l����j��r����^��c1���m6;����|���u����o�[-+��r���|��k��M�s9.�[��K���d)�u:=�W���U*5��v�M&���V�E�q8��_/�K���d�i4�}���_/�K%���Z���a�x.7�������M��y�~��g��l+
��I����V�B ���L#���B�@��P���I�r��F�@  ��\'��B���H"1,��}���o7��f�I$2���G#�H�b�d��t��K%�i�z�g���V�E"1�l�����n�K%�T
%�i���n�K���d����M&3�L�c�X�f��d)*5�V�E"1�l+���b�H"�X�f��d�T
%�i�z��G#���I�r��F�A 0�|�o��m6�].7#�H�b�H���\'��d)*���f�I$�y<����?���q8�������~��g3������X���i4:=������_/�E��x��W���U*��M&3��F��`��T
��I���l+��E�q8<>?���q8<���o7���S���E��x�w����k5�V!��T�e�y<>?�O'����I�r�L���x��W+��r�L#�d����b���B���������@  0��^�G#���B  �x.�[-+
��I���l���z�N�A��X��y����w��n�E��x.���v�c1��V�B�@  �x.�[-�k5�m���~���s��N���p��V��b���B��������@ ��X����t-�k5��v��h�j�e29.��m6�].��m6;������f�I$29.7���a����G���T
���d��t�V��b�d�i�z'�����d)�j�J��A���L����J���`(4:=����z�g3���|�o7�F�`(4�}�����?�O'	"�X�f	��Q(�z�N����X�f��d)��z�N  ��\��s���G#��D���X���|�o�[�V�a�x���}>���w;�N�A�p�v�M��y�~�O����Z����J�B  0�|��w��n��p���K%�T
%����b�d)��z�N�C�P�d�T
�R���A�p,���~��a�x�n�K%�T
�R���A 0�|�o7#�H�b�d��J!�h�j
%���Z�Q(4�}�?���s�\'�D!(4:��O'��d�T
�R�D���D��p�l��j
%�T�����V�B ��X��S��J�a0��^��c1,��}���o7�F ���L#���B��@  �x�����z�N  0��^�C!��T
�����I$�y�~�O'�I��������Y,6��n���X�s�\��s9����~�@���H��Q(4�������}��?�C!���M&3�L��q���O'���R	"�X��S)�j�J�B�@ �p��[-��j�e�y<���_/��e��|�o���v��f�I$29�w;����Z����J��A 08�~����y<>?����y�~�O��i4:=��w;��G�Q(4���_/�K��I$29���}�����o�[�����Y����v��f	��x��W+�e29�n��e29.����[��K��I�r��y<>?�O'	�b������e29�n��b�H���h�u:��O'	������E"1��V�E"�����a0��^�@������A 08���o7�c1,�{�^�C!(4:�^�A�p,��}���_/��b��R�D!(4:�^���q8<����w���W+�������J�P�r���C��H��Q(4:=/�K��I���l�k5-�k�Z�c���F��`��������T����l��u:�^��a��\'�I$�y����w�]�����_/��e2���G#�H"�����a0��^��c�����a08<>?�O'	�b�H����T
���d�i4�}��_/�K%�T�e�y<>?��g3&3����a08�~�O'��B���@�`�h�u����o�[-��u�}�?�A���L#$�y�~��g�Y��[���e��|�o�[��K��I����V!�h�u:=/��������A �x��{��O'��d���Z����p�v��C!��T
��I��Y,6�].�[���e�y<����o7#��R	���h*5-��j�����h�����W+
�R	�b�d�i���n�K%�����f����`(4�����������w;��G#���B�����@���H��x.���v�F���@�`�h�j�J�B  ������q8<��_/�B��P��R�D�����F��`��T
%)*5-+
��I��Y,6;�S)�u:�^���p�v�M&�Y��[���e�y�~�C!�h*��M&��l������W�U*5����m6;�g3�����p��V�E"�X��S)����U*5�m������w;�N�`������i4:�^�C��H"1�l�k��M&3��S)���j�J�����H�b�H�b�H"1���K%�������i�����k5��K���d�i�z����|/���Q(�z�g3�L�c�X&���V�E����������N�C�����A 0���O'	���h*5���[���e���^���p��V�B  0��^�C!(�z��G#$�y<>���w;��s�\��s��N�A���L��q��^��c��L#$29.7����i��].�[-+�J��H��x���k�Z�Q(��].7��f����I$2��N����X�s�\'��B  �x��W�U��z�����M&���V�E��x����u:�^����D�a08<>?���s9.�[���e��|�����~�G���T��r��S�T
%�T
�R�D!����f�I$�y�~�����L���x�����z��G���T
�R�D���X�s9�n�E"�X&�Y,����_/��A�p�l�U*5��v�F��`��Z#�����`�t��v����i4:�^�A �x���}>?�O'	�b���l�k5�m6;����q�|�o7�M&��l+
%��t�m6;�N�C!���J���`(����W+
%)�j��r���C��H"�X&3�f���R���A�p�v��f��d)��U���].7��C!��T
�R��B �p���K%�i4:=�o7�M��y<>?��c�X��y��_/�K%)*�Z����p���K%��t��v�M&3�L�����N��`(4���_���u������{�^�G#��������D�P�d)����U*5��K��I$�y<>?��g3�f��d����b��Y,6;'�I���l+�J�B ��X&3�s��N  ��\��i���n�K��I$2�\�S�T�e��������|��w�]�w;'�I��Y��[�V��b�H�b��D�a08�~�G#���I$2����c�X&3&3��S)��U*5�m��}>����{=/��e29.����[��K%�T�e�y<>?��a�����c1���K����R�D�P�d)*5����m�{=��������w������������z�g3�s9�n������J���D��H�b���B���������H"�X��y�~������^�C!�h�u�}>�_/��b�H���h���j�J��p��V�����������T
�R	�q�|�W+�e29.�[�V�E�q�����s9�n�B��@��P$2���G�Q�t�m���~�O'	��Q(�z��G#$�y<����o���v#��D�a�x���k5�m�{�^����x��W+���b��D�a�x�n��e������s���G��h��U���]�����_/�K�R	"�X������M��y<>��o7�Q�t���[�V��b��R����`��T
�R	�q�|�o�[-�U*5-+�J!�h*5-��u:=�o7�c���F�@  0�|��k�Z�F��P���I��Y,��}�?��g3���C��H���h�����W+��r�L#�d�i���n�K%)���]��{��O'��d)*�����i4��~���q��^�G�Q��Z���a�x�w��n�K��I�r�L�c1�v��C!(4�}�����o7��f�I$29��{�^����x�n�E"��L��q�|/���r&���V!�t��K%��t�������m6;��s��N�@�`�h*�Z����p��V��p���K�R�D!�h��U�u���_��k��M&�Y,6;����|�W�U*5���[-����j�J��H�b�H�b�d���E��x����u:=�o�[�V��A �x���}�?�O'�I�������r�f	�b�r��F�@  08����w����k�Z��C!��T��r�L#$��|�o7�M��y����w;����q8<��������_�W�U���].7��f��B���@  0�|�o7��C�P�����R	���\�S)*��M&3�L�c�X&3��S����b��R�D��p,6�].�[�V����h�u���_���u��~�A 0��^�G#��R��B ���L�Q(�z���y<>?�G#��Y���m�{=�o7�M&3�f���R���A �x�w�]�w;���y<��?�C�P$2��N�`�h�j��r�L�c�X�f	�����J�����A��X&3�f��d��t�m6���W+��E"�X���|/��e�y<>���w;�����^�G�Q(4:�^��a��\'��B�@��P$29���k5�V�B��P�r��S)�u�}>����{��O�S)�����j
�R	�b�d�i4:���g3�L#�H��Q(4�}>���w��n�E"1�v�M&�Y,6;'�I�r��F��P���I�r���������C��H�q8<��?��c��L��h�j�J�B ��X&3�f��d)*5�m6��n���Q���M&��l��u���_�W���U�u�}>?����y��_/�E��x�n��e�y����w������z�N�A �x�n�B ��X��S�T
%�i�z���c��L�c1�l��u:=�o��m��}��_��k��M��y<�����_��k5�m6���W�U*5��v�F�`(4���_�W�U*5-+�e2������x���k�Z�F��P�d�T
�R�D!����E����N�@��P�����R�D����B ��X&�Y,6;���t���[-��u�}>?�O'����I���l+
�R���A 0�|����}�?��g�Y,�{��O'	���h��z�g3�L#������I$2��N�C�P�d�i�z�g����K�R���A�p�l�k5���e2����c��L��q8<>�_��k5-��u��~�O�S)*���f���R�D!��T�e��|��w;��i4:��O��i4�}��_/!(��]���}>�_�W+�J�����H"����C!�t�V�E���\���t-�U*5-���z��G�Q(������u:=�o��m�{��O'	������c1�v#���B�@���H"��L����\'	�q����g��l�U�u:=/�K��I$�y<>?�����|/���r&��l�k�Z���x�w���W+�J�����H"��L������b$��|�W��j�e���^�C!�h�j���b����V��H�b��D��p,�{=�o7�M&�����e29.�[�V�E��x�����z����q8��_�W+�J�P����V�B ��X�s9��W+���b$2�\�g3�L#����A��X����^��c1���K�R��B�@������A����F��P�d�T
%����b�H�q������y��������_/�����T
��I$29�w;�N��@�`��Z#$�y���o7����p���K%�i4�}�?�G���T��r�L�Q(�z�N�����L#�H"1�v���x.7�F ���L�c1�l��j����l�U*�Z�����X���i4��~�O'�I�r��S)�u�}����_�W��j�e�y<>?�A 0��^�G��h�j�J�B���H��x�n��e29��W�U*5-�U��z�N�C���D�a0���O'��d�T
%)�u�}��?�O��i��]�w;��s��N�C!(4�}���?�O'���R��B�@ �p�l�k����S�T
%���E�����G�������Q���M&3&�Y,��}>?���s9.�[-�U*5�m6��n��A�p�l+
%)�����W+����l���z��G#���l��u�}�?�G#�����R�������D�P���l�U*5�m6����k���f��B �p�l+���Y�v�F�@��P����d�T
�R	�q8<��?�O��i�z��i4:=���{�^��P$���^�A�p��[��K%�i�z�N��`���J��A 0�|�W�U*�Z��C!�h�u:�^��c1�l�U*��M��y�~��a0��^�A�p�l�k�Z������G�Q(�z'��d����M&�Y�v����i4�}>������~�C������`�h*��M&�Y����v���T���Y�v�M&3�L�Q(���n�K�R���A 08<���?�G#�����R	"1�l������j��r�f	��Q(4��~���s�\���y�����{��O�S��J����P$�����g�Y�v��f��d�i4:���g3�����p���K�R�D�P�r��S)*���f�I$29�n���r����t�m�{�^�C�P���I�r�s���G�Q�t-�U*5�m6;'	����T�e2��N��a������q8��_�W+�J�������a08��_��k�Z#�d���Z��q��^��c1,��}��_/�a���N�C�P�d���Z�c�X���|�o����[-�k5-�k����S�T
��I���l���z'�I�r��F�@���H��Q�t�m�{���g3��S)�j����Q(�z���c�X�f�D���X��y<����w��n�K%�i4:=���u:=/��b��D�a�x�w;�g�Y,6�]�w�����u:=�o�[��K�R�D!�����b�H�q8��_�W+�e�y<������?�O��i�z'�D!����E"1,�{=�o7�F��@����D�a���N����X&3�s9�w��n���Q�t-+��r&3��F�A 0�|�W+�����h��U*5����m6�]��{=/�B��@  ����G��h�j���b�d��t���[�V!�h�u��~���q8�~�O��i�z��G#�r�f	���h��U*�Z�c�X��S�T�e29�n��b�H����T�e�y��_/��b��D�a����G#���B�����@ �����C�P$29��{�^�G�Q(4�}>���w;'�D!����f�D���X����^�G#�r�����Z�F�@����D�a0��^��c���F ��X���i4��~�O'��B�@  08�~���s�\���y���o��m�{�^�C!�h��U*���f�D�a���N ���L����\���t�m6;��G����J�a0�|/�B��P���I$�y<>?���s��N��a��\'�������D�a08����w;�g���V!���J!�h��U*�Z�c�X&����K�R�D�P�d��J���X����t-���z�g���V��H�b�r��S�T��r���C!�t���[-+�J��A ��\��s���G#���B�`(���n�a0�|���u:=�o��m6;�N�C!(4�}>���w;�N��P���l�U���].7�M��y<�?���q�|����}���������������_/���X�������s����c�X���|�o�[�V�a�x�n�K%�i���n��b��D!��������T
%�T
%)���j����l��u:=����}>?������^�G#��D��H���\���t���e29�n����B�����@ ��X��y��_/�K��I���l�k5-+��r����t�m���~��c1,�{=���{��O�S)��U*5�V����h�u:�^�G#��R����`�h�u:=��w;���t�m6�]��{=/�K�R	"�X&3&��l�k�����i4���_/��e2��N�C��H�b��D�����A�p����v��f�I$��|���{=�o�[��K%�T
%�T
�R���A ��\�g3�L���x.7����i�z��s�����q8<>�_���u����o7���S�T�e���^��c�X�s�\�g��l���U��z�g3���C��H�b���B����@�`�h*5��v�M&3����a�x��{�^�C�����A 08<��?�O�S)�u:�^��c1�l+����l��u�}������{�^��@ ���L#$���^��`�h�������j��E"1�l���z��i4��~�G�Q(4:�^�A�p�l�k5��v����\��s9���}>?�O�S�T
���d)�u:=�o7�Q(��]��{=���{=�o�[-�U*5-��j�e29���}>?�G#��D�P$�����g3�L�Q��Z��h��z�N��a0��^�G�Q���M���|/�K%)��U*5�m�{=/�B���H�b�H�q8<����?�O'����I�r���C��H�b��D!(4:=��w;����|�W��j
%)��U*5��K�R	"�X�s9�w���W+���b��D���X�f����`��T��r&3�s�\�g3�f	�q8�~��@  ��\'	�b��D����L��q��^�@�`�h�j��E"��L��h�u�����w�].�[-+��E"�X��S)�j�J���X����t�m���~�O'�I�r�L�Q(4:��O�S)�����W�U�u��~�C���D!�����b�H"���F  �x������].7��C�P�r�f�I$2�\��s9��W+�J���`��T�e2���G#�d������h�j�J��A 08�����{��O��i����W��j���b�d)*�����i�z�N��P�r�L��q8�����{�^��c�X��S)*��M�s��N�A 08<���_/���Q�����S)��U�u�}>���w���W�U*5�m��������}>��o7�F����@ �p,6����k�Z#$2�����q�|��w;'�D�����A �x����u:�������^  �x�n��b$����O'�I�r���i��].�������[-�k�Z��q�|��k�Z�F�A�p�l�k�Z�F��`(4�����w�����u:=�o�[-��j��r&3��F�A 08��_/����P�d)*5�m6�].7��h*5��K%�i��]��{=/���Q��Z�F��������@ ��X�f�I$2�\'����I�r��S�T��r&�Y��[-��u:=�����~�C!(4��~��g3��F������B�@ ����F����H"1,6;������f	"1��[-��u:����s9��{�^���q�|�o���v�����t���e�y<������{�^���q��^�G��h��U*5����m��}���o7��f�I���l+�J�B��@  ��\'�I$2��N��a�x.�[�����Y,����_/!(4:=/��b$����O�������S�T
�R���A���L#��R	"1�l�k�Z�F�A��X�f	"1��V���`�h�j��r��y��_��k5����m�{=�o7�F������@  ����G#�r�L��q�|���{�^���q���O'�D���X�s���G#�����R	��Q(�z��G#���B�@��P�r�L���T
%��J!������i����W+��E���\�g��l+��r�L�Q(4:�^���q��^�G�Q(��]�w;�N�C!����E"�X&�Y�v���S)�j��r����a��\�S������h*�Z�F��@��P$29�����_�W��j�J��A���L����\'���R	"1,�{���g3�L�Q(4�}����w��n����B  ��\'��d)�j
%��J�B  ���N�C!�t-������W+�J���`��Z�F  08<>�_�W�U*5��v�M�s�\���y��_�W+����Q��Z#��R�D���X���|/��A�p,6;�����x.7�M&3�L��q��^���p�v#�H"1��V��b����d)��z'���R�D!��T
%�����f�D�P���������I����V���Q(�z��G#��Y�v�c1���m6;�����x.�[�V�B ��X�f	��Q(4�}���_/�K��I$�y�~���q���O�S������h��U�u��~��P�����R���A�p���K%�i4:�^�G�Q��Z#�H��Q�t�m6���W+��E"�X�s���G��������h���j��E"�X���i���n���Q(4�}�?��c�X����t�m6;��s9�����_�W��j�e��|�o7�F�@ ��X���|�W�U���]�����_�W+�e29��W�U*5����r��y<>�_/���r�L#�H�b�H�����J�a��\��s�\���y<����_/�a��\'�I$��|����}����w�].7���a0���O'�D����B ��X�f	�q��^���p������Y,6;�N��`(��].�[�V����L�c��L�Q��Z�c�X�f	��Q(4:=����}>?�G#������P�d�T�e2���G��h*5�V���Q��Z��q�|�o���v�M&�Y�v#$29.���v��f	���h��z�N �p��V���`�t��v��f	���h�j��E"��L�c�X�s9����~���s�\���y�~���p����e�y<�?�O��i4:�^���p�l+��E����N��`(�z����|/���D��H�q�|��w��n�E"1�l�U��z���c1�v�������������F�A 08�~��c1��V�E�q8<>���w��n��b�d���Z�����N�C!(���n�K�R	��Q������i4:�^���P$2��N�@��P�r�f�D�P��R���A�p�l+�J!(���n����Y��[-+�J���`��T��r��F�A���L����J�B ��������X�f	�b�d��J��H�q��^��c1�l+��r���C��H"1��V�E�q8<>�_/�E"1�v�M�s9.���v���a����G��h�����j�����h����U��z�S�T
%�i��]�w������z'	���h�����j�������J������D�����F��@ �p,6�]�w���W��j�J��A 08<>�_��k5�V�B��P�r�L#���B�`�h�u:�^�G#�H��Q��Z#�r��F�`�h�j�J!��Z�c1�l�k5������l�k5�m6��n��b���B��@ �p,�{=��w;�N��@ ��X��S�T
�R	�q�|��w�����u��~�A 08<����w;�N  08�����{������|�o���v#�d)*��M�s��N��a��\�g3���C�P��R	���h*��M���|���u�}>?�O'	��Q�t���[����r�L�Q�t�V���X&3���i�z��i�z���c��L��h�j���Y�v�F�@��P$29��W��j
%�i��].7��C!(4�}��_���u:��O'���R	���\��s9.7�c�X&3����t�V�E�q8�~��g3��y<����o7��f�I$2�\'�I$�y��_�W+�J�a0��^��a08�~�G����J�B ������a0���O'	�q�|�W+�J�B�`(4:=�o7���S)��U*����S������h�����j�e2����c�X���i�z�g3�s9��W+�J�B ������a���N �p��V���Q(��].���v�Q��Z����p�l��u���_���u:=/!��T�e��|�o�����m6�����u:=����z����|/��b����V�a�x.7�M&3��F ���L#��D���D�P��R	�q8<>�_/���r�����p�v��f��d�T�e2����c1�l�U�u�}���_�W�U*���f��d�T
%�i4:�^���p�v�F�A��X�f������H"��L�Q����f�I�r��y�~�O�S��J���X�s9.��m6���W+��E�q������y<>��o��m�{=/���r&3��F�@�`����E��x.7�M&�Y,6;���t���[-����]�w;�S)��U*�Z#�H�b��R	��x.�[-+�J������D�a0�|/���`(4:���g3�L#����A�p,���~�O'�D��p�l�k5�V�E"1�v��f�D!(4:=��w;���c�X&����K�R����`��Z�F��@  08��_/�E�q8���������o7��q��^��`���M��y�~��g���V��b���B �p�����r��F��@�`(�z�N ��X�f�I�r&��l�k5�m6��n��e�y�~��g3���i�z�g�Y,�{=�o��m6���W+������T
%)�u��~��c1���K���d��t��v�����t��v#�H�b�H�b�������d�i�z��s9�n����Y�v#��R���A�����C�P$�y<��?�C���D�P��������R�����P�d��J�a��\'	�����J���X�f�I$���^�C�����A�p�v#����d)*5-����]�w�]��{��O'���R	�q���O'�I��Y��[-�U*5�����v�M�s9�n�K��I��Y,�{=�W��j�J!�t�m6;�N  ���N�`(�z�N�C�P����������V����h��z��G�Q(���n�K%)��z�N�@  �x��{=�o7��C!�h�j
%�i��]�w�]����~��c1,��}>�_�W�U�u:=�o�������[�V��A�p�v�F�`(�z������\�g3&3�L��q�|/�E��x.7�M�s�\��i4��~�`����E��x�n��e29�n�K%)�u�}>�����}����_�W���U*������t��v���a08<>����{�^�C�����A �x��{���g3�s9��{��O�S)�u:��O'�I�r��F��������P���I�r&3��F�`(�z�S���E"�X�f�I�r&3��F���P��R��B��@�`����E���\�S)���].7��f��d�i4:=�o7�Q����f	����T�������e2��N�C�P$�y�~���s�\'��B�����@�`�t�V��H�q�|��k5-+
��I$29��W+
%)*5���e29.�[��K%�T��r��F  ��������\�g���V�E"����C!��T
%)��z������O'�I$29�n��b���l+�����h*���f	��Q(4��~��g3�L����\�g3�L�c���F��@�����B���H�b$�y<>�_/�B��@ ��X�s���G�Q�t�m�{=��w;�N�A�����C!�h*��������M���|���{=�����].�[-���z��i�z��G#�H"1���m6�].�[-+
��I$29.7�F������A ��\��s9.�[-���z��G��h*5���e29�n��b�H�b���l�k����S)�j
%�T
����R�D�a0���O��i4:�^����x���k�Z�Q����f	�b����d)�j
%�i4:��O'	������c�X��S�T�e��|�W�U*5�V������D!�t����m����_�W+�J�P��R	��Q�t����m��}�������w��n�E"1�l�U*�Z��C!�h��U��z�N�A ��\�g3���i���n���Q(�z'����I$�y<>?���q8<��?���s���G�Q(4:=�o���v�M&3�f��d)*5��K��I$�y<>�_�W��j
%���Z�F�@ ��X�f�I$�y<�����o�����m�{=/��p,�{=/������C���D!(��].7��f	������E"1,��}��?  0�|��w�����u:=��w;'�I�r����t-�U��z��������i4�}>��o7����i�������z����Z��C!(4�}����_��k5�m6;�g��l+
�R	�b�d��t�m���~��g��l����].7�F���@ �p�l�U������k5�m����_���u:�^�C��H"����C���D�a���N��@���H�b��D!(�z��G#�d��t�m6�].��m6;'	��Q�t���[-��j�e2�\����Z����\�g3�L���x�n�B �p,6;'�I$��|��w�]���}>�_�W+����Q(4�}����w;�N���p���m��}�����{=/�K���d�T
��I��Y,����_/�������P�r�L#�d)�j����Q��Z�F��@ �p�v��f�I$2��N���@�`�h��U*��M������g3�s9��{=��w;�S)��U�����W��j��E"1�v����p�����[�V���D��p�v����J�B��@�`�h�j�J��A���L��h�u��~��g�Y,6�]��{=�W+
�R�D�a���N��@�`���J���X&3�����O'�I$�y<�?���s��N�@ ����F ���L��h��U���������].��m�����o�[�V�E"1�l�k5���[���e�y<>����{=��w�]�����_/�K%�i4�}>?�O�S�T
�R���A 08<�?�`����E�q8�~�O�S)�j
%����M��y<>?��g3������M�s9��W�U�u�}���������o�[��K�R	��Q�t��K���d�i4:=��w;���y��_�W�U�u:=�o�[�V�a�x���������k�����i�z��s�\������O�S)�j�e2�\'��d����b�H�b�d��t�m6;�N�C!(4��~�O'	"1�l����].7�c��L���T
%�i4�}>�_�W+�J��p�v�c�X�f	��Q(4�}>������~�������O'��B  �x��W+�J�a�x.7#�H�b�H��x��{��O'�D������C!�����b��D!���M&�����e29.7�F�@  0��^�@  0�����s�\'	����T�e����O�S)������k5�����Y��[-�U*�Z�F���P��Y,6;'�I���l��j����Q���M&�Y,6;�����^�����\�g3���C!�t�m��}��_/��b�H��Q�t-�k��M���|/�a0��^�G#��D!�h��U*��M����^��c���F������A�p���K%)�j��E�����G�Q��Z#$2�\'�I$��|�o7�M��y<��_/�K%)*��M&3�L���x.7�M&�Y�v��h�j��E"1,�{=�o7��C����B  �x�n��A ������q�|�o�[�V���Q(�����k������t�V�E��x��W���U����n��e2�\��s�\'�I�r��F�@��P$2���G#$���^��a0���O�S)���]�w��n�E"�X&3���i4:���g3��F �p�l�k5��v�Q(��].7��C!�h�u�}>���w;'�I$���^����D!��T
%�T
%��t�m���~�G#�H"������p�l+����l+��E������c1��[-��u:�^��c1�����r�f��d��J!��T����l�k��M���|�o7���S)�j�J�B�`(4���_/�B��@  �x���k5-+����l+
%)���j
%)�u:=�o7���a0��^�G�Q�t������[�V�������E"��L#�������H�b$2���G�Q(�z����q��^�G�Q(�z�S)�j��r���|�W�U�u��~��g���V���Q(���n���r&��l�����U*��M�s��N���p�v��C�P$29.��m6��n�������K���d)�j
%���Z�F  0����g3��F�`�t���[�V��A���L��h�j
%��t��K�R	����T
%�T
%��t�m�{�^��c1�l��j�e�y<������}>?���q8�~�����L#�r&3��F��`��T
�R	�b�H����N��a���N  ����G#�H��Q�t-�k�Z��C�P$2�\�g��l��u�}>?��g�Y�v�Q��Z�F����@�`���J��A 0�|/�K%�i4:�^���P�r�����O'���R�D�P�r�s�\�g�Y,6;�N�@�`�h����U*5��v��C!�h*5�V�E�q8�����{�^����X&3�����p�l��j��E"��L#���B  0�|/�E"�X��y�~�����L#��������Y,�{��O�S�T��r�L�c1,��}>?�A �x��W�U��z�N�C�P$2�\�g��l+
%�T
%�i4�}>��o�[��K���d�T
��I�r���C!(�����k�Z���a08��_�W��j�e�y�~�O'	�b����A ��\�S)��z������f���R�D�a�x.7�M��y�~���s���������G�Q(�z�g3�s9.�[�V��A���L���x��{=�o7���a08�~��`�h�����j
%)*�Z���a��\���y<���������{�^�A�p�v�M�s������x������]���}��������_/�����l��u��~�@ ����F�`����E"�X�s9�n��b�H"�X�f�I��Y,6;�����x.�[����r��y��_/����Y���m�{=�o7�M��y<�?�`���J!��T
%)�j�����h��U*�Z����p,��}>?���H�b$�����g��l��u:��O'�D����B���@ �p�v�M�s9�n�E"1���K%)*5-����j������T�e2��N��������a��\'	�q8����w;�N�����D!�h*5�m�{=/�B����@�`(4��~�G#$��|��w���������W+����Q�t-+���Y,��}�?���q8�~����y<>��o7�M�s9�n������D!���J��A 08<�?�O'�D��p�l��j��E�����G#��R	�q8<����w�]��{�^�G#�H�q�|�o�[-+�e�y<���������_/�B����@ ��X�f	"1���m��}�?�O���t�m��}������������w�]�����_/�E"1��V�E�q�|/�K%��t�m6�].��m6;���t���[-�U*�Z��C!�h���]���}���o7��f	"1,6�]���}��?�G�Q���M&3�f	"����C�P��Y,6;�N���@��P$29��W+
���d��t-���z��G#$29�n���D��p�v����i�z'�I�r��F��`��Z����p�l�������k5��K%��t�m6��n�K���d��J!��T�e�y��_��k�Z�F��P�r�������L�����N�@  �x�n��e29�n�K�R�D!����E��x�n��A�p,���~��g3��S�T�e2��N�A��X�f����I�r�L��q8<�����_�W�U*5-�k��M��y<>�_���u�}>?�O'�D!��T��r����t���e29�n��e�y�~������F��P�d)*�Z��C��H�b$29��W�U�u:�����y<�?���s9����u:=��w;'��d)*���f�������������I�r����a08�~��g3��S)*5-+
��I$29.7����i4�}>���w;'	���\��s�\�g���V���X�f���R�D��H"1,6;��G��h*�Z��C���D��p��V�E"1���K�R�D!�h*�Z�c1�l+
%)��U*�Z�F  08<����w��n�K�R	�q8���o�����m�{=��w��n�K%��t��v�F����H�q�|/��e29���k5-+
%���Z��C�P����d���Z�����N�C�P�r���C!(�z��G�Q�t�m6�].7������Z�c1���m�{�^��c�X&3���C!��T��r��F�`��T
%���E"�X�f	���\��s�\'�I$2�\�S��J�a��\��s��N�A 08�~��g3&3��F��`���������M�s9�n���r��������y<>�_���u�}>����{��O���t�m6;�����^��a�x�n�K%)*�Z��q�|���u:=��w;����q8�~��c1��V�E"�����a08<���_/��e��|��w�].7�F����@��P$������s��N ���L#�����`����E�q�|/�K%�i4�}>?�G#������P�d���Z����p�l+
%��J�B��P$�y��_��k�Z#�H����T���Y����v#$��|�o��������m6���W��j
��I$�y<��_/�B�@ ��X������M&3�f��d�i4��~�C�P�d�T�������e��|�o7��f��B �p,�{=���u�}���_��k5�m�������{�^���p�v����p����v��h��U*5�V�E��x��{=�����~�G�Q��Z�F��@ �p�v�F�A�p,��}��?�C!�h*�Z#����A �x�n!(4��~�G#����d��J�a08<��?�A ���N�`��T����l�U�u���_�W+�J!(��]��{=/�K���d���Z�c�X�s��N�C!�h�j��E"�X&�������Y�v����p��V�E�q8<��?�����������\'���A �x�w;�S)�u�}���o���v�M&3�L��h��U*�Z��q8�~����X�f�D�a����G��h��z�����x�w��n��b��Y�v��q8<�?�G#�r&��l�U*5��K%��t��v��f�I$29.�[���e�y���o7�F��P�d����b���I������e29����u��~���q8<>?���s9�n�K%��t��v��f��d��J����P�r&��l�k5�V�a�x.7�M��y<��?�G#�H���h��U*�Z��C!���J�P����d��J�B  ����G#��R�D!(4:�^�C!(�z����q���O'����I��Y,���~����H�q��^��`�h�j��E"��L���T
���d��t�V��H�q8<����o�[-�U���]�w�].7���x�n�K%�i4:�^���@������A��X���|�o7��f��B�`(���n���Q(���n��e�y�~��c�X����t�m�{�^���q8�~���s�\�g�Y�v�M�s9�w�].7�M&3��F�`��Z��C!�h��z�N��`�h�u��~����y�~�O'��B�@  ����G�Q���M&�Y,�{��O�S)*�Z��C!(4��~�O'	�����G�������Q��Z����p������Y,�����o�[�V��b��D�P��R��B�`�h���j�J���`�h*���f	�b��D!(����W�U��z��s�������\�S)���]���}>?����x.����[���e����O����Z�c�X��S����b�H"1,6�].��m�{=�W�U*��M��y<�������?���s9�w�����u��~�O'��B���@�`�t-�U�u:��O'��B�@�`����f�I$����O�S)��U*5���[-+�������J�B���@���H��Q(���n��b�r�L����\�g3�L#�r�����p,�{�^�G#$�����g3��F�A��X�s�\'����`�h�j�e���^�C�P$29�w���W�U�u:=�o������v��C!�t����r�L���T�e29�n��b$2�\��i4:=�W���U*5��K%�����f�D����L�����N����X��������S)�j
%��J�a08����w�]�w���W����j
%�T���Y�������v�M��y<>?��g3���|/��e�y�~�G#�H�q���O'	�b���l�k�������Z�����X�f�I��Y��[-+���b�H��Q���M&�Y,�{������|�W�U�u:�^���p,�{��O�S�T�e2���G#��D�P$����O'����I��Y,��}���_/�E"��L���x�n��A �x.7���S���E����N�C!�h*�Z�c1�v�F�����D����B���@ �p�l�����n���������Q�t�m6���W+
�R�D�P�r��S)*5�m�{�^�G#�H��Q(4��~�C!����f	"1���K�R	��Q����f��B�@  ����G#�H�q����g��l�U*�Z�c��L�������c�X�f��d����b�H�����J���`���J��A 08<�?�O'����`��T���Y�v�M����^��c���F��`��Z�c1�v��q��^�C�P$29���k5�m���~�O'�I���l����]�w������z'	�b��D!(4:=���u:��O��i�z'�D��H"��L���x�w����k�Z�c1���m�{=���{=���u�}>���w����k��M���|/�K��I$�y<>�_���������u�}>?���q��^�@  08<>?�@���H�q�|�o7��C!(4:=�W+������T
���d�T
%��t��v#�H"1,6��n��b�����`(��].7�c1,���~��c���F�`��Z��C!(��]���}����_�����]�w;�N�C!��Z#�H���h�j���b��Y���m��}>�_��k5��v��f	���\'��d�T
%�i��].��m�{=/�K%�i4�}���_/�K%)����U��z���c��L#����d��t��K%����b$��|/�����F�@  08<����_/�K%)����U*5�m6����k5-�k���f�D�a0�|�o��m�{=��k�����i��].�[-���z��G�Q(�z���c1�l���z�N��a0�|�W���U*5��v�M�s9�n�B ��X&3��S)���j
%��t�m6;���y<>?�O�S��J�P��R	�q8����w;�S������h*5��K%�i�z'��d���Z�F��`�t�m�{�^����D!(���n�B ������a08<��?�C��H"�X&3�f�I�r��S�T
%)*5�m���~�����|/����Y���m�{=/��b�H�b�d�i4:=�W+
�R�D�a�����c���F ��X�f	�b���B��P$29�w���W+��r��y<��?�G#$�y�~��c1�l��j�����h�u:=���{=/�K%��t-��j��r�L�c1�l+�J�a�x�n�E�q��^�`��T
�R	�����G�����E�q8�~�C!(4����o7�M��y�~�C���D���X&���V����L�������c1�l���z�������g3���|/�P$�y�����{=�o7�M�s9.�[�����Y,��}���o�[-���U�u��~��c�X�f���A 0�|�o�[����r�L�Q(���n��e��|�o��m6�]���}>�����}>?��g3��S���E�q�|�o��m����_�W+�J��p�v�c��L�Q�t-����]��������{=�o�[����r�f������R	�����J���X��S��J!�t���e29��W�U*5��v�F��`�h�j�e�y�~�O'	"�X&3�L���x.7�F�`��T��r�L�Q(4����o�[-�k5-�k5-�k5�V��p,�{=�o����[�����Y,�{�����y<>�_/�E�q8��_/���`���J!�t��v���S���E�������q���O'�D!�h�j���������Y�v�F���@�`�t���[���e�y�~������F�A 0����g3�L�Q(�����k�Z�c1���K%������S��J���`���M&�Y��[-���z��i4�}>���w�]��{=�o��m6��n�E"��L�Q���M&�Y,6;�N����X&��l+���Y,6;���y�~�@��P$2�\'	"1,�{�������^��c��������L��h�j�J��A�p�l�k5�V�B���H"�X�����Z�F�@ �p���K%�i4:=/���Q(�z���c����C������`����f	�q8<�?���P$���^�������C��H���\�g�Y,6;�N�A�p�����r����a�x���k5�m���~��g3&��l+�J�P�r&3�s�\������f�I��Y,��}>?�O'��d��J����P�d����M�������s�\�g�Y,���~��g3��y<>?���s9��������{=�W+�����h��U�u:=��w�].7�M�s�������\��s�\'����I���l+��������E����N�C!(����W�U����n�B��@�����B��P��Y,��}>?�O�S)*5�������m�����o��m6;'	�q�|�o�[�V������J��p��V����P$29��W�U*��M&�Y��[�����Y,6�]����~����y�~�`�h*5��K�R�D�a0�|�o7�����t��v���S���E"��L�c�X��y<�?��c�X��y��_/�B������@  ��\'������R	�q8��_��k5�m6;��s�\�S)�u�}�? �����C����B��P$2��N������@ �p��[��K%�i�z��G#�d)�u�}>��o���v��q�|�W�U*5��K%��t�m�{�^��`�t-���z'����I$2���G#�H"1�l���U�u�}>��o���v�M��y<>?�C�P���������I�r��F�`�h�j��E"1����v�c���F�A ��\�g3�f�I$29���}>?��`�h��U��z�S)*�Z����J�P�r���i4:=�o7���S)�u:����s����c������p,6;'	��x��W�U*5���[-�k5��v��C��H���\�g3�s9��{=�W+�J�B ��X&3�L�Q�t�V�E������c���F��@�`(���n��b�d�i�z�N��a0�|�o7��h�j
�R	�b�H�b���l+�J��A��X�f	���h*�Z�����X&���V�P��R	�q�|/����Y,��}�?���@��P����d���E��x�n���r�f�I���l�U��z��G�Q�t��v�M&�����e2�\��s9�n�K�R�D�a���N�C!�t-��u��~�C���D�a���N�C���D�P$2�\��i4:=��w;��G#��Y��[��K%��t��v�F�A���L#��������D�a08�~�C!��T
%���Z��C!����f	"1���m6��n��e2��N��@�`�t�����v�F�����D!(4:=�o�����m6��n���Q���M���|��k5-�k5�V�E����N�C!�t�m�{�����y�~�O'	�q8<>?���P�����K��I$�y<>��o����[��K�R�D�a��\'�I$���^�����\���y<>�_����z���y�~���p�v�c1,�{�^��c1�����r���C��H���h��U*5�m�{��O'������R�D!��T
%��t����m�{=���{��O'	����N��@��P$���^�C!(4:�^�C�P��R�D�a0��^��a�x.��m6��n��b�H�����J���������`�t����������m���~������A �x.7�M���|�W+���b�r��F�����D��p�l�k�Z�F�A�p��V��b��D��p���K�R��B����@�`��T����l�U*�Z�Q�t�m�{=�W��j��r��S)���]���}���o�[-��j����Q(������u�}�?��g�Y��[-�������U�u�}>��o7�M��y������}>���w;�N����H�q�|���u:=�o���v�F���P��R	�������q8<��?�O'	���h��z��i4:�^�C!�h*5���[�V�B  08�~�G#�H"1��V�E�q�|�o7�c1,6;�����x�n��A�p������Y��[��K�R����`����f�I�r�f�I�r�����p�l+���b��R�D!���M&3&3�L��q8��_/�B�@���H���h�j�e2���G�Q(����W��j
�R	�b�H�q8�~��g3���i�����k5�m6;����|/�B�@  08��_/�K%)���j�e29����~�G#�r�L��h*5���[�V�B��@  �x�����z��i��].7����p,�{=�o���v�M��y<�?���q8�~�O'���A�p��[-+��r�f����I$���^�G#���I�r���C��H�b�H��Q(�z����q�|��k�Z�F�A��X&3��F�����@�`(�z��G#�H���h��U*�Z��q�|�o7��C�P�d��������t�m6�]���}��?����y��_/�����l��u:�^ ���L�Q���M&��l��u����o7��f�I$�y�~�O'�����P��R���A �x��{����s�\�g3�f�D��H�b��D!��Z��C���D!�h�j��E"1�l+
%���Z�c�X���|�W�U*���f�I�r&��l����j��E�q8�~�G#$2���G#���l��u����o�[-���z�N�@  �x�w;�g3&3�f�I��Y,6;�N  ��\�S)*5�m6;�N��a0�|��k��M�s�\�S�T
�����I���l+���b�H"1,��}�?�O��i4�}�������_�W����j�e2�\�S)�u��~��a0�|�o7�M&3&���V�E"1,�����o7���T
�R�D����B�@��P��R�D�a�x��{=/������J�B�`��Z�Q(��]�w�].���v�M&3�L��q8��_/�K%���E"�X��S)�u:=�W+�J������������`�t�������V�E"1�l�k��M���|���{�^�C!�t�m6;�N�C!�h�u:=�o7#�H�b�H��Q(4:=/�B�`��Z�Q(�z��s9�n�����l��u:=/�K%�i4:=���{��O�S�T
���d����M�����O��i4���_/������`��Z��q8���o7������Z����p���m����_�W+�J�B �p�v�M���|�o�[�V��A��X&3������X�f	"1�v�c�X&3�L��q8<���o7�F�@ �p,6;�g�Y,�{�^�G�Q����f	�q8<���o�[��K%�i4:=�o7��f	"1����v�F�A��X&����K%)�j�e���^��a0�|/�K�R	�b���B�@  �x.7#$��|/���r��F��`��Z�F���P���I$�y�~�C�P$�����g3���|�o7��q��^�A���L����\�S)���j�e2�\����|�W+
���d���E���\��i�z����|��w;'��d��������t�V�E"1�l+�J��A�p�v�M&3�f��B���H��Q(4:�^�@ �p�l���z�g3����a��\�g3���i�z����q8�~�G��h��z'����I���l�k5�m�{�^�C!�h*5��K%�i���n��e�y<>?����@�`�h*�Z�F���@���H�b�H��Q(4�}>?�C��H����N�A 0��^�`(��]�w;'��B �p��V�E"�X�f�I$�y<��?��g�Y,�{����s9����~��c���F��@��P��R�D�a08�~�C��H��Q(���������n�E�q8����w;��i4:=�W�U*�Z�F �����C!����E�q8<>�_/�B�@����D��p,�����o7��f�I�r�L#��R��B ���L�Q���M�s��N���p�v��f�����P�r����a��\���t�m�{=�o���v��f	"1,6;�N��a0��^ ����F�@�`�t�m6�].7�M&��l+�e29.7��q������y<�?���q�|�o7�������F��`���J!��Z�F���P�d)�j�J�a0�|�o��m���~�O����Z���x.7�M���|�W+�����V�E"1�l��u:�^�C!�t-��j��E���\�S)����U��z�N��a08�~��g3�����p���K�R	���h*5��K�R	��Q(������u:=/�K%����b��D!��Z��C�P�d�������T
�R	�����J�B�@ ��X���i4:=/���X�f�D!��T
%�i4����o7#��D��H��Q(�z���t�����Y���m��}���_/���r��S��J��A 0�|/�K%���E�q��^�@  ��\'�I�r�L#�d���Z�c��L#�r��F���H����T
��I$����O'�I��Y�v#�H"�����a0���O'�I$29��{=/����h*�Z�Q(�z�N�C�P�r�L�c1�v��f�D�a�x�n�K�����I$�y<��_���u���_/��e2����c1���m6;��G��h*5�m6;�S��J!(����W+�e�y<>����{��O'���A �x�n�K�R	�b�H����N��a��\���y<����_/������D�P�d)��z'�I$�y<�?�O�S)�j��E�q�|��w;�g3��F��`(���n�K%�����f	"�X&�Y�v�M��y�~�G��h���j�J!��Z�F�@ �p���K�R�D�a�x�n���Q(�����k���f�D!(�z�������g�����e��|�o7��f����I�r�L�Q��Z��q8��_/��e�y�~�G�Q(4:�^���q���O�S�T���Y,��}>���w��n�E�q8<>?�O'�I�r���C�P�d�i4:=�������W�U*�Z��C!(�z����q�|��w�����u�}>��o7�c��L#�H���\�g�Y,�{�^�G�Q(4��~�O'�I$2�\���t�����v��C!���M���|/����Y��[-��j�e�������y��_/�K�R��B  �x��{=/��e�y<>?�G���T��r�f�D�a�����c1��V�E��x.�[��K%)���].�[��������K%)�j�J�a0���O'�D!�t-�k5�V�E"����C�P$���^�G#�H������c1��V�B�@��P�d��t�V���X�f��d�i4:=��w�]������o7���a08��_/���D�P�d��J���X�s�\��s9���k5-����].�[�V��b�H"1�l+��E��x.��m�{=�W��j�J!�h�j
�R	�q8���o7��f�I�r�����Z#�d)�j
%�i4�}��?�C��H�b����d�T
%�i4:=��k5��v��f�D����B�@  ����G�Q(4�}��������?�O��i4:���g�Y,6�].���v��f	"��L�Q(�z�N�A 0��^�G�Q(��]��{�^��c���F���@ �p�v�M&�Y����v��f�I�r��S��J�B  �x.7�F  ��\'����I$2���G#�d)��U��z��G�Q(���n�B����@  0�|/�B�@ ��X&���V�����T�e�y�~�O'��B ����F�@  ���N���p�v��f�I$��|�o�������[���e��|����}>�_/�E�����G#�r���i4:=�o7��q8<>?�O'������H�q8<>?�O�S����b�d)�j
%�i���n����h*5��K%�T�e��|�W�U�u�}>�_/�K�R�����P�d)�j��r&3&�Y�v�c1���K%��J��p��V��p�l�U��z�N��P����d��t��v�M�s�\�g���V!���������M�s9��W��j
����R�����P�d��t��v�F�A��X����t��K�R	��x.��m�{=/��p�����r��S��J�B ��X�f�I$�y��_/�B�@�`�h*5�m�����o�[-��u:=�o7��f	��Q(4�����w�].�[��K%)�j�e�y<�����_�W�U*��M&�Y�v#��D�a0��^���@�`�t��K����R�D�a�x.����[��K�R��B����@ �p,6;��G#���B�@�`���M���|�o7�Q�t�V�E"�X&3�f�D!��T
�R	"1��[-+�e2�\'�I$����O'����`�h*��M���|����}�?��g3�f	��x�n���`�����S�����Q����f�D��p����v#�H��Q(�z��G�Q���M�����O��i4��~�O'	"���F�A 0��^��c1�v#�d��t����r���i4�}>?�O'��d�T
%)�u�}�?��g�Y,�{�^�G#�H�b��D�a��\�S���E"1�l��u:���g3���C�P�d)���]�w�]�w;��G#�d)�u:=�����~�������A 0��^�G#�d�i4:=/����h*5��v����\���t�m6��n���r�L�c1,6;��G�Q�t���[�V���Q��Z����p��[��K%�����f���R	���h�j�e�y<>?�O'��B��@ �p�l+���b�d��J�a��\�S)*5��v�F�`�h�j�e���^�C��H���\'	"1����e�y������}���_/�K�R���A 0��^�G���T�e29�n�B ���L#�����K%��t��������K%�T
��I$�y<>�_/�������K%�T
�R�D�a0��^�G������b�H�b�H"�X���i4:=����}�?�O��i����W�U����n���Q(�z'	���\'��d)��U�u:����s��N��P��R	"��L#�H�q���O'��d)���].�[-�k5��K%��t������[����r���C�P�r�L�c��L���x�n�E"1�����[��K%�i������u:=��w;���y<���������?����x�w�]�w�����u:=������_/���r����^���p,6�].�[-��u���_�W+�J�B��@  0��^�G���T
%)�j�e2��N���P��R����`����E"��L#�d�i���n��e29�n���Q��Z�c1�l+�e2���G�Q����f���R�D�P$�y���o�����m6;��s9�n������J����L#�H�b��R	�����G�Q(4�}>���w;�N�C��H��Q��Z���x�n����h��z��G#��D!�h*5�����v��C!(�z��G�Q�t�m6;���c1,�{=�W+�J��A�p,6�]��{���g����K���d���Z�F�A 0���O'�I$�y�~�O��i4��~��c��L������G#�����R�D��H�b���I$29�n��b����A 08�~�G�Q�t�m�{=�W�U�u�}�����w�]��{=�W+�e�y<>�����}>�_���u:=/����h*5��K%)���j�J��A��X&�Y,����_���u:=�����~���s�\'�I$29.7��h�j��r�f	"���F��P�d�i4��~����y<�����_/�K�R	"1�l���z'	��Q(�z�N�@�`���M��y<>?������B �p�v����p,6�]�����_/�B��@ �����C�P����d�i4:=/�P$�y��_/�����T�e29���}>?���s9�w;'���R	�q8������}>���w;�N��@ �p�l���z��s���G�Q(����W+�e��|/�K�R	��Q(�z�N���p,��}>��o�[�V�E��x.���v�Q(4�}>�_/��b��Y�v�M��y<��_/��b�d�i4:�^�G�Q(�z�N  0�|�W+
��I�r�L#��D�a��\�S)*5�m�{=/���r�����p�l+
���d����b�r��F��`�h*�Z#��D�P���I�r��F��`����f�I$29.7�F�`�h�j
�R	������c���F �p����e2��N�C��H��x�w�]��{=�W�U�u�}>�����}>�_�W��������j��E�q�|��w;�N�C�P���l��j
��I�r��F�@  08<>?�G�Q��Z�Q(��].7�F�@���H���\�g3�s��N��a�x�w;��s9���k�Z���a��\���y����w;����q���O�S)�j�e2�\��s�\�S)�����j���b�r��S)�����j
%)*�Z��C���D��p��[�����Y,6;�N��a08��_�W��j
%)���].���v��f	�b��D�a08<���_��k5��v�F�A ����G��h�j�J����L�c����C��H���h��U�u�}���_�W+��E"���F�@�`��T
%��t��K%)��U*5-�U�u�}>�_����z�g����K�R	�b�H�b����d���E�q������y<>?�O��i�z��G#��D�a�x���}������?��g�Y,�{=�o7�c1,�{��O�S)��z'��d�i��].7�F�����@�`(����W+
���d�T��r���i�z'���R	�q�|�o�[-�U*��M&�Y�v����i�z�N�A����F���H���h�u�����w�]���}>���w;�N��`���J!��Z���T
%)�j�J��p�l�U���].�[���e29.7����p����e2������x�n�������K%����M�s9.�[-��u:����s9�w;'��d)��U*5���[-�k5-�k�Z��h*5��v��C����B��P�d�T
%)*�������Z�c1���K%)�j
��I$29���k�Z���T
%�i�z���y�����{�^��P�r�f��B �p�l����].��m�{���g3��F����@��P������e�y<>���w���W�U*���f�I�r����t-���z��G�Q(�z'���R���A 0�|��w���W�U*��M�s�\'��d)�u:=��w;�g�Y,�{�^�C!���M�s9.��m�{������|�W��j�e������s��N�A 08��_�����]��{=��w��n��e�y<>?���q�|/�K%)*����S)�j���Y,�{�^�A 08��_����z��G��h�j�J�P$2�\�g����K%��t-+��E�q8<���?���P�d)�u���_/��e2�����q8<>?�O'�D�P��R�D!������i��].7�����X&���V�a�x��W�U*5-�k��M&�Y,6;��G�Q��Z�F����H"�X�s�\�g3&�Y����v����i�z�g3�f�����d���Z��C��H�b�H��Q��Z�c1,�����o�[�V!(4�}���?��g3��S)��z�g��l+��r����t�m6��n�K%�i�z�N��a��\�g3���C!�h*��M&��l�k���f�I$2����c1��V!�h��U*��M&���V�E"�X��S���E�q8<�?��g3&3�L#�d)�j�e�y��_/���`(4:=����z�S���E��x����~�C!�t�m���~�G#�r����a�x�n�K���d��t��v�F��`(�z'	�b�������d�i4����o�[�V!�h��U*���f�D���D��p�l+���b�H�b�H��Q�t����m��}>?��c�X�f���R	"1,6��n�����H��x��W�U*��������M&3��F  �����c�X�f��B�����@ �p���K��I�r�s���G����J!�h�j�e29.�����m6;�N��`�t�m����_/������J�B�@ �p,6����k5��K%�T
%�i4:=���{=��w;��s��N�C�P$���^ �p�l+��E����N��P$��|�W��j
%�i4:=�o�[��K%�T
�R	��x�n�E"1�l+���b��D��p,6�����u������{�^���q8�~�O�S����b$����O'���A�p�v����\�g�Y�v���S�T�e2�\'�I���l+�J�B�@��P����d�i����W+�J�B  08�~��c�X�f	�b�H�b�d�i���n�K�R��B  ����G�Q(4��~�O������f	���\�g�Y������m6�]��{��O�S�T
%�i4:=/�E�q8�~�O'�I��Y�v����p�l���z����|�o7�F �p��[�V��p���m�{�^�����L#�H���h������U�u:=�o7�F ��X��S�T�e��|�W+�J��p�l+�e��|��k�Z����p,6�].7���S)��U*�Z�c���F���P�d�i4�����w��n�K%)��U*5�V�E"1�l�k5-��j
���d�T
%����M�s9�n��H"�X&�Y,�{����s���������G�Q(��].7��f	���h��U��z���c���F��@�`�t-�k5��v�c1�v��f�D�a�x.7��f	��x�w���W��j��E��x�n�B��P$2���G�Q����������f	�q8<>?��g��l�k5���[-��u�}>?����y�����{�^��c�X���i��].�[��K�R�D�a�x��W+
���d�i�z�g�Y�v�����t���[-��u:=/����h*�����i��]�w���W���U*��M&�����e�y<>?�O'	�b���l�k5��v�F�@��P$29�����_/�K%)�u:����s�\�g3&3��F��`�t-��u�}��_/���`(��]���}�?�G#�d�i4�������}>���w;'�I$2�\�g����K��I��Y�v�F���H�b�H���\'��d�i��].7�F�A 0�|/�K%��t-�U��z�g3�L���x.7�M&3�L#�H�b��R��B�@����D��p�v��f	��Q(��].�[��K��I�r�L����\�S)*5�V��b�������H�b�r�s�\'	"���F �p��[��K%�i4���_��k��M&�Y,���������~���s9�w;����Z�F��`���J�a�x��W+
%�T
%)*�Z#���B�`����E"1��[��K�R�D��p��V���Q(�z�N���p,6;�g�Y,������w�].���v�M&3��F���P�����R����`�t���e2�\��i��]�w��n�K�R	�b�H�b�H"��L����������J��A �x.7��q��^���H���\�g�Y�v�M&���V�����T
%)*��M��y�~�O'�I$2�\�g3�s�\�g3�s9����u�}��?��g3��F��`��T���Y�v��h*5��v��f����I����V�E�q����g�Y����v��f	�q�|�W��j�e2�\'��d)�j�e2�\�S��J�B��@ �p���K�R�D�P�d��t-��u��~�G#�H"��L�c1���K%)*��M�s9.7����p�l�k��M�s9�������n�E"�X&��l��u:�^���p�v�M&3����t�����v�����t-��u��~��c�X&��l��j���b�d���Z�c��L���x.7��C!(��].�[-�k5�m�����o7��f	�q8���o7�F  08<����?�G�Q(��]�w;�N��@ �p��[�V�B�������`��T�e2����c1��V��A 0�|����}������?�G#���B ��X��S)*5-�k5���e��|��w�].�[-�U�u���_/�B�@�`�h�j������������T
%�i�z�����x�n�K%)*��M&3�L#�H�b����A����F��P���I�r�L#��D����L���T��r��F�`�h�j�������J!���J!��T
%�i������u:�^����X��S�T
������d�T�������e�y<>��o���v�M&3�L��q8<>?��g3�L�c��L#�H�q�|/��b��Y,�{=�o7�M�s��N��a��\��s9.7�M&3��y�~����X�s�\'	���h�j�����h*�Z#��Y,6�].��m6;'	���h����U*�Z�F��`�h*5�V����L��h�j
%)��������U�u:=/�����A��X�f��d�T
%�i���n�E"1�l��u:��O'	"���������F��@��P���������I�r�f���A�    T          P                                           ��������    �������  �                                  �����������       �����������       �����������       �����������       �����������       �����������       �����������       �����������        �yw        ��   �       L       ��L���x�w�].��m6�].7�F���H"�X�����Z��C!�h�j�J����L�c1�l+�e���^�G��h���].�[����r��S�T
�R�����P��Y���m6;�����^���p��V������D�P��Y,��}��_��������k����S�T��r���C!�h���j��E"1����v�M&3��y�~����y���o�[-+�J����L�c��L������G�Q(�z��    �N���@  �x��W+�e�y�~��a�x.�[-+��E�q�|����}����o7�M&3��F �p,6;����|�W+����l��j
%��J��A���L#�H�b�H"1,6;���t�m�{�^���P�d�i��]����~��a�x�n��e2�\�g3��y<>�_�W��j��E���\���y�~�C��H��Q(�z�g3&3�L�c1,6;��G#�������H�b���I$�y�~��c�X�s9���k��M��y<>���w;���c1�v�F�@���H�������q8�~��g3����a0�|/�B�@ ��X�f	�b���I����V�B��@ �p,6���W+
����R	�����J�a�x��W+
���d�i4�}>?�O��i�z'	���\�g���V�E�q8��_/�������K%���E"����C�P�d)����U*5���e2�\�������g�Y��[-�����n���`(4:�^���p�l���U�u:=�����~�O'�D���X�s9�n�K%�i��].�[�����Y����v�����X&3�L#��D�P�d���Z����J��A�p�l�������k5�m6�����u��~��`��Z�F�@�`(�z��i4�}�?��c�X&3�f����`�h��z��s9�w;'�I������e�y<>?�G#���I$���^�G#��R�D�P$�������y��_/�K%���Z#�H�b�H�����G#��D��p��V�E"1�l���U*5����r&�Y�v�M&���V�E"��L#$2�\�S��J��A��X&�Y�v�M�s9��{�^���q��^�G#$�y<>?���q��^�G#�H��x���}����w;��G#�H�b$2�����q8<���?�O��i4��~�C!���M&3��F���P$�y<����������w��n����Y,6�������].��m�{���g3�L���x���k5-+
�R	��Q���M��y�~���s����c1��V��b����V����P�r���i4:=�o��m�{=/���r�f	�����G�Q���M&3�L�Q�t���[-+�J����B��@ �p,6;���y�~�G�����E�q8<>?��g3��F��`��Z���x.��m�{��O'�D��p,�{=�W+�����h*�Z��C!��T
�R�D�a�x������o���v#�d�i4�}>���w����k5�V��A�p,6;��G#��D�a�x��{=/���Q(�z������O'�I$2����c1,6��n��p,��}>?�G��h��z�S�T�e29.�[-+���b$���^�A�p�v�F  �x�n�K�R	�b��Y�v�M�s9��W����j��E"1�l�k5�V���Q(4:=/�B����D�a�x��W���U*���f�D�a0�|��w������z�N�C!(���n�a��\�S)���]�w���W+
�R�D�a���N���p�v�F��`��Z�F�@�`(4:=����z�N��P�d)�j
%����M��y�~��g���V�B  08����w���W+�J�B�@�`��T
%��t�m��������}�?�A���L�Q(�z�N�C�P����������������d��J!�t���e��|�W+�J�B �p��V����B ��X�f�D���X&���V����B�`�h*���f	"���F���@ �p�v��f	����N�A�p�l���z�N�@�`��Z�Q(4�}�?���s9������o���v�M&3������X�s9��W�U�u�����w;���y�~�G�Q�t�m6;���c1�l��u��~��g�Y�v�c�X&3�L��q8�~�O�S����b�H��Q�t���e2�\��i4:=�o7��C!�h��U�u:=�W�U*5-�k�Z�c�X�s���G#��D�����F�A ��\'�I�r�����p�l+��E"1������������Y�v��q�|/�B  0��^�C!�t�V�B ��X�f��d��J��H"1�l�k�Z�F��`���J!(���n����P��Y�v��C!�h�u:=/�K%��t�V��A 08<>��o�[-+��r�L#���B  08���o������v�M�s�\��s9.��m��}>?�����|�W�U*�Z#�H�q�|/��A 0�|��w;�N��a����G�����E"1�v�����X��S�T�e�y��_/�K��I$29�n��e��|�������o��m6��n!�t����r���i4:=���{��O�S�T�e2�\�S�T��r�L��h���]���}>�_�W+���b����������d��J��A 0��^�G�Q��Z��q����g�Y,�{�^��c1�l�k5�V�E"�X�s9.7�����t-�k�Z��C!�h��z�N�C!�t�V��A��X�f�I$��|�o�[-��u�}>��o����[�V�B��@ ������a�x����u�����w�]�������w;'��d�i4:=��w;����|��w��n�a0�|�W�U����n��e2�\'�D!�h���j
%����M&3�f��d�i4:��O'�I�r���C!�h�j�J!��T
%�i�z�N�C���D���D!���M&3���i����W�U*���f�������D!(���n�a�����c1�����r���C!�h��U����n��e2�\���y�~��c1��V��b�H"1�l�k5����m6�].����[-�k5-�k��M&�Y,�{=���u:=�W�U�u�}���������_��k5�������m�{=/�E�����G��h�u:=�����~���p�l��j�J�a��������\�g��l�k��M&3�s�\���t����m�{�^��c�X�s���G#��Y,����_���u:���g����K�R	�q���O'	���\'���A��X����^����X&3����a�x�w;�N��a08<��?�����|��w�����u��~�O'�D��p,6;��G��h*��M&�Y,6;'�D��p,�{���g�Y,6;�S�T
%)�j�J�B �p�v��f��d)�u:�^����x��{=/�B  0��^�C�P�d�T
%��t��v�Q(�z��������G#�H���h*�Z��C��H"1,�{=/���r�f�I������e2�\��s�\�S)��U�u�}>�_/�B��@  0��^��a�x.7�F�@�`��T
%)�j��E���\���y�~��g�Y,�{�^��c1���K�R����`�h�j
��I�r�L��h�j�J�a0��^�����\�S)*5-���z�g�Y,6���W+�e29���k5�m6�������].7�M&��l�U*5���[���e2�\'��d���E����N����H�q�|��w�]�w�].7#�d)�j�e2�\��s�\�g3�L��q8�~���P�d���E"��L��q��^�G#�d���Z��C!�h���j
%�T���Y,����_��k5-+�J���X����t�m6�].7�F��`��Z��h��U�u���_/�K%���E"1�l+
%�i��]�w;�g3&�Y,6;�N�C!�h�j����Q�t�m6��n�E����N��`��T
%�T
%)��U*�Z#�H�b��Y��[��K%�����f	�b��Y,�{�^�A������a�x�n��b�������r���i����W+��E"�����a0���O�S�T
%)����U*�Z���a����G�Q�t-�U�u:�^�A 08<>��o7���S)������U�u��~��c��L�c�X��y��_/�E"1���K�����I$�y<���_��������k5-�k5�V��p����e2�\����|/�������B�@ �p���K���d�T
%�T
%���Z�c1��V�B �p�v�����t-+�J�B�@�`�h��z�N����H��Q(�����k5�m6�].7�M���|�o��m�{�^��a�����c1�������v�Q��Z���T
%�i4:�^����x.7�F�@��P$��|/��e2���������G��h�j
%)�j�����h��U����n��A 0��^�G��h�j
�R	�b�H�q8�~�O'	�����J��p,���~�����|�o��m6��n�B���H�b��D���D�a0��^�`���J�B����D���X��y<��?��c�����a��\���y<>?���q�|��w;��G#�����`��Z��h�����j�J!�h�u:=/�E"�X&3�f���A�p�l��u�}>������~�O'�����d�i�z�g�Y,����_��k�����i4:=�o�[-���U*��M�s�\���y<>���w;'���R�����P��Y�v����i4�}>����{���g3&3��y<���_��k�Z�Q�t-�k5�m�{=��w;'�I$29��W����j�J��A�p�l���z�N��`����f	"1�v���S)�u�}��?����x�w�].7�F�`�t-�k5�V����P$�y�~�O'���R	�b�r��y<>?����x.���v�F�@���H"������p�l��u:=�W�U*5���e2�\'	"�X�s�����q�|��w���W��j��E"1�l�k5�m6;����|/���`�h�u������{=�o�[-�k5�V��H���h�j�e�y<>?��g3����^  �x�n�K%����b$�y<>?�G#��D��p,��}��?���p�l��u:=/�K%�T���Y�v��f��d)�j����l���z�g3���i4�}���_����z'�I$2�\�g�Y�v���x��W+�e�����g�Y�v�F��`�h������k��M&����K����R��B���@  �x���k5��K%�����f���R	�b���l+�J�B �p�v��h�j�J�a����G#�����`�t-+�e29.7�M�s9��W�U�u:=���{�^���q8<���_��k5-�k5-+����Q(�z'�I����V��b��R	��Q(4:���g3�f���R�D�a��\�g���V��A��X�f��d�i4�}�?�O��i�����������k�Z��q��^�`��Z���a���N�@  �x����~��`����E"��L�c�X���i�z�N���p�l+�e29���k5�V��A �x�w�].7���x������o7�M&3��y<>?�O'�I�r�s�\�g��l��j
�R	"1�l����].��m�{=��w����k��M��y<����_/�K%����M����^���p��V���X��S)�u����o�[-+�J�P$��|�o7����p���K%)�j�J�a08���o�[-�k5����m��}���o7�F�`(4���_/�������K%�i�z�N�`�h��U���].7��q�|/�a�x�n�K%�i4:=�o��m�{��O'�I$2��N��`�h�j
��I���l����].7��q����g3&3��F�@�`(�z��G��h��U*5�V����B��P��Y�������v����i4�����w��n�B�@ �p�v�F�A�p�l�U*�Z�c1�l+�e��|�o���v��f���R	����N��@ ��X&����K�R	�b�d���E�q�|�W+���Y,��}>�_��k5�m��}������?��c��L�Q(�z��i��������]��{�^��a0���O�S�T��r�L�c���F�A 08�~���p,6;�N�����L#�d��J��p�l��j�����h*5�m�{����s��N���P��R	�q8�����{=�o7���S)�u��~�����|��w��n��e��|�o7���S��J��H�b���B�@�`��T�e�y�~��g�Y,�{=��k5-�k5�m6��n��p,6�].�[���e2�\���t��v�M&���V�E"�X�s�\�g�Y,6;'	"�X�f�I$�y<������w�����u�}>�_/�E"�X��S)���j�J!���M&��l+
��I$29.7�F��`�h�j�����V��p���K�R�D�a�x�n�K��I�r�L�����N�C!�h���j�J�P�d���Z���T�e�y<���o�[�V��A��X�f��d��t��v�M����^����X�f�I�r���C�P$29���}���������o�[-��u:��O'��B��@���H�b$2��N�C�P��R��B�@�`�����b$��|/���r�L���������T�e2��N�C���D��H�b�H�b$�y<>?  08�~�G���T
%�i����W+�J�����H�q8<>?�O�����M���|��k�Z�F��@�`(4�}��������w;���y<>�_��k5���[�������V�E"�X&�Y����v��f�I����V�B ����F ����F�A �x.�[��K��I�r���i4���_/�E"1�l���z'�D�a��\�g3��S��J���`���J�P�d)��z�S����b�H"������p��[-+�J�B�`�h���j�J�B�`�t-�k�Z����\�S�T
��I�����K%)�u�}����o�[�V����h����U*���f��B�@�`�h*��M�s��N��`�t�V�a�x.�[�V��H�b���B�@ �p,6��n��e��|�o7��f	"1,�����o��m6���W+�J�B�@  �x��W��j���b����A �x.7����i4��~��g�Y,��}>��o�[-�k���f��d)������k5-���U�u��~����X�f�I�r���i�z�g3��S�T
�R	"����C!��Z#�H��x.���v��h��U*5�m6;��G#��D���X��S)*5�m6�].�[�V���Q(4:=�����~�O���t�m6;���y���o�[-�k��M&����K�R�D������C��H�b�H"1��������V�E�����G#�r&3�f��d��t-�k5��v�F ��X�f���R����`��T
�R	"1�l�U��z'�I�r&�����e�y�~��g�Y��[-�k5�V�a0��^���p��V��A�p�����[-+��E"�X�f�I��Y,6;��������G�Q(���n��b��R����`(�z����|�o�����m��}>?���p�l�U*5-���z�S�T
%��J�����H���h*5-�k���f�D������`�h�j�e����O'�I$��|�o7�F�A�p�l����j���b���I�������r��y<>?�@����D�a�x.7��q8<�?��g3�L#���B�@ ���L�c���F��P�r&3��F�A�p��V��b�H��Q(4��~��`�h�j���Y,6��n�a0�������|/�K%��t�V��H�b$2����c��L��q8��_���u��~�O'�����P$2�\���y<���?�O���t�m����_/�K�R����`����f	���\���y<��?�G�Q(�z���c�X��S�T
%�����f��d�i��]��{�^��a08��_���u���_������n���D�a0�|���u�}>���w;��������G�Q��Z�F�@ �p,��}>?�O'������R�D��p,6;��G��h�j��r�L#�����`(�z�N�C!(4:=/�K�������R	�q��^���q8<>��o�[��K%��J��H�q8�~�G��h*5�m6�]���}�?�O'��d����M��y��_��k5�m6�].�[-�k�Z����J�B �����C�P�d)*5�m6;'	�b�H�����G��h�j
%�i4:���g��l����].7�M�s9.�[���e���^���q�|�W�U*5-����].�[����������r��F����D�P����V���Q�t��K%�i4�}��_����z�g�Y,6;��s���G�Q�t-�k���f�I�������r���C!������i�z�����M�s9�n�K%�i4�}�?�O'�I$�y�~�O����Z����p���m6����k��M&�Y,���~��g3��y��_�W+
�R�D�a��\�g3&3���i�����k�Z����p�l+�e29��{=��w;��G���T�e�y<����w�]���}�������o7��f��d���Z���a��\'��d�T
%)�j
%��J��H�q8<�?��g����K�R	"�X�f��B����@�`��T���Y,�{�^��`��T
%)��U*�Z�F�����D!�����S��J��p�����r��y<>?  ����G#���I$2���G�Q(4:�^�G#��R	���h��U��z�g�Y�v��h�����j�J��A���L��q�|/�E"�X�f���A 0�����s9�n���r��S)�j����Q��Z�F�����D�a�x�n��e���^����x�w�]�w�].�[�����Y��[-+��E"1����v��C�������P��Y,�{=���{�^ ��X&3&3&����K�R	�q8<������?�O��i4:�����y���o��m6;�����^��������a0���O'��d�i��].�[-��u:��O�S)�u:=��w;�����^���q8��������_�W+�J���D��p�l����]�w������z�N�C!�h�j���Y,�{=/�B�`�h*5�m6�]�w�].��m��}���o7�F�@  08�~�O'���A�p,�{����s9�n����Y�v������Z��q8<����w;�g�Y���m6��n���r�f��d�i4:�^���P�d�T�e2���G�Q�t��K%)���j��r��S)��z��G#��Y�v�M��y��_/����Y,�{=�o��m6�]��{=�W+��E"�X&�Y��[���e2�\�g�Y,���~�O��i���n��b�H���h*5�m6�����u:=���{���g3�s�\�S�T��r���i��].�[�V��A�p�l+���b����A 0���O�S�T
�R	�b�H�b�H�b�H��Q��Z#�d����M&�Y,6�].7��f�I$29��{�^����X��S)�����j��r�L��h�j��r�f��B�@��P�r���C!��Z�Q��Z��C���D!(��].��m�{�^��`���M&�Y,�{=/�K�R	"1,6;�g3��F�A��X��y<>?�O'��B����@  0�|�o���v�M�s�\�g�Y�v#����V�E��x���}����o7��f�D�P�r��F�A ��\����Z�c1��V!����f	"1���K��I$��|/���r���i4:=�o��m6��n���r��F���@�`�h������k5�m6����k5����r�f�I$29�n�E�q8�~�G#�H�b����V�����T���������Y,6;���������t���[-�U*5-+
%��J�B���@����D���X�s�\���y<>�_/��p,6;'�D�a��\��s9����u:=����}����?����x�n�K�R�D��H��Q(4:�^����H"1,6;���c1�l+�J�B��P�d���Z��q�|��w;�N���P���I�r�L#�H�q�|�o����[-�k5�V�B�@��P����d�i����W����j�J�P���I$��|/����P�r�L#�d��J��������H"��L#�����R�D!���J�B��@  08��_/��b$2��������N�����D!���M&3�����p��V�B�@��P�d�T
��I������e2��N���@  0���O'�I����V��A 0�|��k5�V�E�q8��_�W�U*5���[-��j�J�a���N�C!(4����o��m6;�g3��F ����F��`(�z�N��@  �x��W+�J��������A��X&3��F�A 08<����w;��i�z�N��@��P���I$���^���p,6���W���U�u:��O'���R���A 0���O'��B�`��Z��C!�t��v�F�`�h��U*5���e�y�~��g3�L����\������O'���R�D��������p,6;�N�C�P�r��F  08�����{=�o7����������i4�}��_/��e2��N�C�P�d���E"�X�s�\�S)���].�[�V�E"1���K%��t-�k5����m6;��i��].7�M&��l��j�J��A 0�|/�K�R	"1,�{���g3���i�������z��G�Q����f�D!�t������[-+�J��A 0�|�W+
%�i�z�S)�j�J����P�d)��z�N��`�h��z��G#�d��t�m6;�N ��X����t��v��f��d�i4����o�[-�k5-�����n���Q(4���_����z'��d�i4�}>��o7�F�@�`�h����n���Q(��].7��f	"1�l�k�Z��C!(4:=����}>?�`(4:�^�A 0����g��l+�e29�n���`�����S�����Q�t�m6;�N����X���|��w;�S����b�H��x�n�����l+��E�q�|�o��m�{�^���p�l�U*5�m�{�^�C�P�d�i4:=�W+�e29.7�c1,6�].7����i4��~�O��i4:�^���p�������v�M&3�f	��Q�t��v��q8���o7�M�s9.�[�V�B �p���K����R	�b$2�\�g3��F  ��\�g�Y,���������~�G#$�y���o��m�{=�o����[-�k��M&3�L�c�����a0�|����z����q��^��c1,��}�?�O�S)*5��K��I��Y,�{��O'�I$29.���v�M&3���C�P����d�i4�}>��o7�����t-��j
�R��B����@�`�h�j������K%�T���Y,6;���y<����?������^�A�p�l�U*�Z��C!�t����m6��n�E"��L���x�n�E"1,6��n�E"1���K%�T
�R�D�a�x��W+��E"1���m�{���g3�L�c1,6;��G�Q(4:���g�Y���m��}�?�G�Q�t���[�V�E"1��V���X�s�\�g3�L#��D�P$2��N�A ��\��i���n����Y�v��q8<>��o7����\�g3�s9.7�Q(4��~�O�S��J�B ���L#�H"���F�A�p�l+��E"1�l+�J�a��\�S)��z�������N����X&3��S��J��A �x��W+��E"1,��}>?���@�`(�z��G#�H�b���l����].�����m6;�S)�u:=/�K%�i4�����w;���y����w;'�I$2�\'�D!�t���[-+
��I$�y���o7����p����e2���G#��R	�b����d���Z�F�@�`��Z�c1������Y�v�M&3�L�c�X�f�I$�y��_/�E"1��V�a08<>?�O�S)�u:=/�a�x���k5���[-�U*���f��d����M&3��y<��?��c�X����t�V�B�`����E��x�n�K%)�j��r�s�\�S�T
%)*5��v�F���@  08<��_/��e�y<�?  08�~�@ ������a0�|�o7�M�s9�n��b�H"�X���i�z'�I$��|��w;������f�I��Y,�{=��w;�N�@�`��Z���x���}>��o7#��D�������a08<��?�G����J��A�p�l+�J�����H"�X�f�I$2���G#�H��Q�������t��v��f	�q8<��_/��e29�����z�N �p�l��u:=/�K��I$�y��_/��e�y<>�_/!��T�e��|/�����A��X���|/�K%�����f�I$29.7�F���P�d)�j��E"���F�@  ��\�g�Y,�����o7��q8�~�C�P�d�i4�}���?��`�h�j
%����M&3���|/!������Q��Z�F�@�`�t-��u�}������o��m6��n!�t�m6;���c�X&3�L#�d�T����l��u:��O'	"��L�Q��Z�F���P$�y<>����{��O�S)�u�}����w;��s9�w;��s9��W�U*5����m6�]��{��O'���������R	�b�H�b��D���X&3�L��h�j�J��p����v��C�������P�������d�i4:=�W�U*5�m6;'�I�r&3���C!�t�V�E"��L�c1�l�k�Z�F��`�t�m6;��G����J!��Z��q8<��_/�K%)���j��r���C!��Z��h*�Z#���I����V������J��A 0�|�o7����p,�����o7����J�a�x���k��M��y<>?����y<����_/���r���C�P�d)�u��~�O�S)���].7���x����~�O�S�T
�R���A 0��^  0�|��k�Z#�r�f	"�X�s9�w��n��p,���~�����|/��e�������y<>����{=��w;��s9.7�c�X�s���G�Q(4:=���{��O'�I����V�a�x�n���r���C!�h�j���b�d)�����j���b�r���i4���_/����h��z'	"1�v�c�X���i4���_/�B�`�����b���I$2�\'�D�P�r���|�o7��f��B�@����D�P���I��Y,6;'�D��p�l�k�Z�F�A �x��{�^���p�v�M�����O'���A�p,�{�^����x�����z�S)�j
%�i��].��m�{�^�G#$29�����z�N�`�h������U��z'�I$���^��c1,6;���t���[-���U�u�}>�_/����Y,6�]�w���W�U*5��v�F���P$��|�W+�J�P��Y,6;'�I�r��y�~�O'�I$2��N  ��\�g3�����O�S)�j
%���Z���x��{���g3&3�L#�H"��L���x.���v�M&�Y�v�M&3�L���T
%��t-+��E"�X���i�z'���R	��Q��Z�F��`�h��U*5�m��}���_/�K�R	���h*��M�s�\������f	"��L�Q�t�m�{=���{=������_/���r���i���n�E"��L�c�X��y�~�O'	�q8<>?�A 08<������?�O��i4�}��? ��X&���V���Q(���n���r���C��H�q��^�G�Q�t�����Y����v�M��y�~�O�S�T
%)�j�J��p��������[-�k5��K�R����`(4���_��k�Z�c����C!(4�}����_/�E�q��^���q8<>�_��k5��K%)��z��G����J�B��@  ��\�g����K%����M�s��N�C!�����S�T
%)���j��E"1�l�U�u:�^�G����J�B�@ �p�l�U�u:���g�Y����v�M�s9�����z�N��`���J��A 08���o�[�V����h��U*5�m6��n��e29�n��������e��|�o7�F���H���h�u:=������_/�E�q�|�W+���b�H"1�l+������T
�R�D���X&3&�Y,6�]��{��O�S�����Q(4:=�o7�F�A�p�l�k5�m��}>?��c1��V�a0��^���p��[-�k��M�s9.�[-�k�Z��h�j�J���X&��l��u�}���?�O�S)*�Z�c��L#$29�n�����T
%�i�z���c�X��S�T
�R	�b����d)*5��v��f�I���l��u:��O'��d�T
%�T�e2��N�`(�z��G#�d�T�����V�E"�X&��l�k�Z�����N�A 08�~�C!�t�m6������z'�I$2������x�n���Q(�������z�S�T
%����M��y�~�O'������R	��Q(4:=�o7����i��]����~�G#���B �p�v��f	��Q(�z���c1����������������e2�\�g3�s9��{����s��N�C!�h�j��r��y��_/�K%���Z�F�A�p�v����\'	�q8<>�_/�K%��J�a�x��W�U�u��~��a��\�g�Y,�����o�[�V���D!��T
��I���l��u:��O�S�T��r�f�D��p��[�V�E"1,6�]�w�].���v����p,6��n�K%�T�e�y<>?��g�Y��[-+�����V�E�q�|����}�?���q8<����?�O��i4:��O��i4�}>�_/�B�@�`�t�������m6;'���R�D����B �p�l�k5�m6��n�����T�e�y<>?���s9��W+
%�i4�}�?�O����Z�F��@  08<>?��g3���C!����E"1�l�U*5��v�����t�m6;��G#��R��B�`��T
��I���l�k�Z�F�A��X�������f	��Q�t��v�c��L���T�e29���}����_/�K%��t��v�M&�Y,���~�G#�H�b�r���C�P�������d�i��]���}>?��g3��S�T
%��J�P�d�i4:=�o7��f���R	�b$�y<��_/�B�`(��������].7#�d�T
%���Z�c�X�f��d)�j
�R	����N���p���K%�i�z�g3�L�c1���K%)�u�}�?��g3�L����\'���A��X�s��N��a�x�w;�S�T
%)�j�J�a�x.�����m�������{=��k����S)��U*�Z��C!�h����n��e2��N�A�p��V���Q�t�m6;�N��@��P$�y���o�[-�k5�V�E�q�|�������o�[-�k���f����I�r�s9.�[-�U��z��s�\���t��K%����M�s�\�g3&�����e�y<>����{��O'	�q8<>?�G#$2��N�C��H�b$2�\�S)�u:=��k5-+
�R�D!�t���[�V�E����N�������@�`(4�}>?�G����J�B �����C!�h���]��{=��w�].7���S)��U�u��~����H"1,6�].�[���e2��N���P�d)�j�J�B��@��P�d�T�e��|���{���g3�L�c������p����v��C!(4:�^�G#��D�a08��_���u:=�o7�M&���V��b�H"�X��S)��U*�Z�F��`��T
%�T
��I$��|��k���f	"1��V�E��x�n�K%��t��K%���Z#�r���i��]��{��O'�I$�y��_/��b$�y<>?��a�x.�[-��u����o7�F��`���J!��Z�c��L��q8�~ �p,�{�^  0�|��w;�S)�����W��j�e29��W�U�u���_�W�U�u:�^�G#�d�i4:=/���r&�Y��[�V!��T
%�T
��I$2���G#�H�b�H"1���K%�i4�}���������o��m6��n�E�q8<>��o�[-���z���y�~�O���t-+������T����l+�e���^�C��H"���F�A��X�s9.7���a��\���y<>�_�W���U*5�m�{�^�G#�H"�X&��l����].�������[-�k�����i4�}>�_/��b���l�k���f��d�i4�}>?�C!�t��v�M�s��N�C!��T����l��u��~��@�`����E���\�S)���].���v��f�I��Y�v�F ��X�����Z�c���F�@ ����F����H���h�j
%�i4:=���u:���g��l+
��I$29��W���U�������u:�^����x����~�C��H��Q���M&3��F�A�p��V�a08��_/�����l����]��{=�o7���S)����U������k��M����^��a08<��_��k5��v�F��P��R��B��@���H�b�H�q��^�G#��D�P����d�i���n�K�R	�b�H�b��R��B�@��P��Y�v����i�����k5-��j���b��Y,�{��O�S)������U��z�N�`(�z�S�T
�R��B�@  ��\��s9�n��e2�\�S)���]��{=�W�U*�Z�F�A��X&3&�Y�v#$29�w;�N��a�x��W+
%)�u�}>?�O'	�b���l��u�}>�_/�K��I�������r�L�c1�l����].���v����i4�}�?�O'�I$29�n�K%)�u���_/����Y�v������Z������L#�d�i��]�w��n���Q�t-�U��z���c�X�s����c1���K%�i4�}>?���P�d����M��y<�?��g3��F����@  0��^��a��\��s��N�C�P�d)�����j
�R	�b�d)*�Z��C!�h���]��{=/��A ����G�Q�t-+����Q(4:=�o7#�H�b$�������y<�?���s��N�C!�����b�����`(4:=��w����k�Z��C!(4�������}>?�O'�I$29��{=����}�����o7�M�s����c1,���~�G#$�y�~�O'	����N�A 0�|�o���v��f�I$�y��_/�K%���E"�X���i����W����j��E�q�|��k5��v�����X��y�������~�@ ��X�f���R�D��H������c����C!����f��B��P�r�f��d��t-��j��E"1���K���d���Z�c���F�A��������X�s9.7���S)�j�e�y<��_/�K%�i��].7��f	��x��W+��E"�X&3���C���D�a0��^���q�|/��b$�y��_/���`�t�m�����o7�c1���K����R�D!(4:=��k�Z���T�e���^��c1���m��}�����?�O���t��v�M���|/�E�q��^�G����J�B �p���m6����k�Z��h��U*5-����]��{���g�Y,6;'���R�D�P�d���Z��h�u�}���_��k�Z����p����e������s9�n���r�f	�b�d�i��]���}>��o�[-+����Q(��]�w;����q���O�����M&3��S�T
�R	"�X����^�����\'��������B  0�|��k5-��u:=�o7#�H"�X&��l����j
��I$2���G#��D!(4���_�W+���Y,6�].����������[-�k�Z���x�w�]�w�].���v���S)*5��������������v��h*5-��j�J�B  08���o��m�{=/����Y�v������Z��C!(�z����|���{=��w�].7�F�A�p�l�k�Z��C�P�r�L#�H�b�H"1�l�k��M��y�~�������O��i��]����~�O'�����d)����U����n��b��D�������a08�~�O'�I$29��W�U�����W+������K%��J����P$2�\'��d��t�V��p�������l�k5�V�E��x.�[-�k��M&��l�k���f���R��B  �x�n���Q�t�V����h�u�}��_/���Q(4�}>?�O'�I�r�f��B����D��H"��L�c��L#���B���@ �p�l��j�J�a0�|�o�[-�U*��M&��l�k5�V��A �x�n�K%��J��A����F�A�p,�{=��k5���[��K�R	�q8<�?�C!(��]�w�]��{=��k5���[-+���b�r�f	���h�j�e�y�~�C!��T
%)��z�N  ���N�C!���J����P�r�f��B �p�v�M�s9.7��f	�b���B������@�`��Z��h������U*��M����^��c���F ��X�s�\'��d���Z�F��P�d�T
�R�D��p�v���S�T
�R��B ��X��S�T����l�k��M�s9.��m6;��G#�H�q8�~�O'�I$2�\�g���V��H������E����N�@  0������y<>���w��n��A 08���o�[����r�L�c1��V���Q�t�m�{�^�A����F���P�d����b��D�a�x����u��~�O'�D!�h��U��z�N��a�x�n��b�d�i4��~�O'��B��P$����O��i�z�N�C!(4��~��g3�L�Q���M��y<>?�O����Z�F�A 08���o�[-��u:=���{=��w�]�w;���y<>?��c����C!�t�m�{��O'�D�a�����c�X�����Z�F����H"1�v�M&3���|�W�U*��M��y��_�W+
%�i���n��e29.��m�{=���u:=���{=/��b���l�����n�E"1�l�k�Z��h�j���b�H�b���B����@����D!���J�B���@�`�h*5���[-��j��r��F ��X���i���n��p�������l�k�Z����\'�I$�y<>����{=�W�����U*5��v��h�u��~�O'�I$�y<>��o7����p�l���z�g�Y,�{=��k���f��d�i4:���g3&�Y���m�{=�W��j������T��r�������L��q8�~�C���D��H��Q(���n��e29.7�c�X���i4:=��k5-��j
%�i�z�N�C�����A����F�A 0�|�����~��g3�L����\��s��N�C!�t�m6�]��{=�W�U��z���c1�v��C�P�r��F����D��H�b�H���h�j��E"�X�f	�b�d�i���n�K%�T
�R	���h�j�J�a08<>?�O�S�T���Y,6;��s��N���p��V���D��p��V�����T�e��|�o������v��f�I$��|��w;�g��l�k�Z�F  0�����s9�n�K%�i�z��G#����d�T�e�y<����w����k5�m����_/�K�R	"�X������g3�L��h*5-�k5�V����P�r�f�I�r���C�P�d��t��K%��t-��u�}>�_/�K��I$��|�o�[���e�y������}>?�G#�H���h*5�m��}>?�O��i4��~������F �p�l�k5����m6;�N����H�q8<���?��c����C�P��Y���m6�].�[���e�y<>�������_/������C!(�z�N�@  �x�w���W����j�J����P�������d)����U*5��v��h�j���b�H��Q(4:=�o��m��}�?����y<����o7�M�s�\�g3�L#��R�D����L�Q(4�}����������o7�M&�Y�v�c�X&3�L#��D!�h�������u��~�����\��i4:�^�C��H�b��Y��[�V�B�@�`�h������U�u:�^�G�Q(4:=�o7��f���A�p�l�U*�Z����p,6;���c�X��S)�u:=�W+��E���\'	"1�l�k5-�k��M�s9�w;�g�Y�v�M���|��w���W�U��z�g���V��A��X����t-�U�u:��O'��B������A������a0���O'	��Q(�z�N����H�q8�~���@�`(4�}��_��k5���[�V�����T��r�������L�Q�t�V�B�@ ��X�f	�q�|/��b$2���G����J�����H�b$��|���u��~�G#�H���h��z��s9.7�c1����v����i4���_������n����B�`����E"1�l�k�Z�c����C!����E��x��{=�o7����p��[���e2�\'��d�i���n��b�H�b��D�a�x�w;�N��a0���O'�����d)��z�N��`�t�m6��n��b�r&��l�k������t����m6;'�I$29����u�}>?���q8���o7��C�P�r�s9.�[-����].�[-+
%�T�e�y��_���u:���g�Y��[��K�R	�b�r�L�Q(�z'	�b��D!�h���].���v�c1,�{��O'�I�r���i��]�w;'�I�r�L�c1�����r�s9��{=���{��O���t���[���e����O�S�T�e�y���o7�M�s9�n�K%����M�s9.7�M&��l+�e2�\'���A�����C!�t-�k5���e2��N�C!�h�j�����h�j�J�B  �x�n��H�����J�B  �x�n���`��T�e�y�~�G�����E"�X�f�I$�y<�?�������G#��D�P�r&�Y����v�M&3�s��N������F���P���I�r��������F�A�p��������V�����T
%�i4:=/�K�R	�b�d�i4������{�^�G#�d�i4��~�O'��d�T
%�i���n!���J!�h�u���_/��e��|�W+�J!�h���j
%�i��].�[�V�E"1�v��f�I����V���`�h��U*5��K%�i4:=��w;��s��N��`(�z'��d)��z'�D!���J�B����@�`��T�e29�w��n�K%����M��y<>��o7�M�s�\��s���G������b��Y�v�F��`(���n�����T�e�y<��_/�E�q8<�?�A�p,6�����u:=����z�N  08��_/!���J��H�q�����s9��W+
%����������M�s��N�C!���M�s���G#�H�q8�~�����\���y���o7�M&3��y�~�����|/��p�l+����l�k5-��u:������|����}>?�O��i�z���y����w���W��j�J���D!�h*5�m6��n��b�H���h���].�[�V��b���I$29.�[-��u�}�������{=�W+���b����V��b����A�p����v�c1�����r���C!(�z�N�@  �x���k5���e2��N�C!(4���_/�������K%)*�Z�c1�l����]�w;�N��@  0�|���{���g�Y,�����o����[��K��I����V�E"1���K�����I�r�����p,6��n��e29.�[��K����R	�b��D���D!���J!��T�e2����c1�l+�J!�h*�Z�F����H�b���I�r���C!���J�a�����c1�v��q8<>?�G#�r�L�Q�t�m�{=����������z�N  08�~��c���F��@�`(�z�N���p�v���������T
%�T��r�������L�c��L#���l��j
�R	�����J���X�f��B  �x.����[��K�������R	�����G#�H��x�n�K��I�r��y<>��o7#$2�����q8<�?��g3���i4:=��w;�N �����C!���J���X�f	��Q(4:�^��a08��_��k�Z���x.�[-��u:=/��e��|��w�]��{�^�A�p�l+�e2�\'�I$2�\�����^�`�h�j
�R�D!�t�m6;��G�Q(��]���}>�_/���������r�s9�w�]�w���W��j�e������s9���k��M�s�����q8<>��o���v��������f����I$2�\��i4:��O'����`�h�u:�^���p����e2��N�@  0�|��k�Z��C��H�q8<>?��g3�L�c1���K��I$2�\�S�T
%)����n��b���I$�y�~�O'�I$�y<����o����[-���z�g��l�k5���[-+�J!�t��v�F�A���L�c1����e2�\��s9�������w��n�K%)*��M����^���p,6�].�[-���z�N�A ����G#��R�D!�h*5-��u�}��?�O����Z��C!(���n��b���l�k5�V�E���\�g�Y�����[���e��|�o�[��K��I�r����a08�����{��O'	�b��D����L���x.7���x���k5-��u:��O'	�q�|�o��m6�]����~�O�S)�u��~��g3������X��y�~��c�X�����Z�c1�l�U*�Z#$�y��_�����].7����i�z������\�g�Y,���~�C!���J��A�p�l��u�}>?�O'�I$�y��_/������C!����f�I��Y�v�M&3��F���P��R�D��p�l+��E"1��V�a��\�g�Y���m�{=������_�W+�J���`��Z#�H�q�������|��w;�g3���|���{�^�G�Q(�z�g�Y�������v��f	����N��a0�|�W+��E"1�l��j��E������c���F �p�l�U�u�����w;���c�X&3�����Z��q8�~�A 08���o�[�V�E"�X&3�L�Q�t�����Y�v�M���|���{=�o�[�V�a0�|�o7��f�D����L�Q(4�}�?����y<>�_��k5�m6�].7���S�T�e�y�����{=�o�[�V!��Z�����N���p,6�].��m6�].7���a��\��s�����q8�~����y�����{=���u:=����}>?��g�Y,�{=�o��m��}>?�G��h���j��E"��L�c1�v��C�P�d�����f�I��Y�v�Q(�z���������y����w;��G#�d�i�z�N����H"1�v�c���F����D!��Z��C����B�@ ��X&3���C!�t���[��K%��t-������������W+��E�q8��_�W��j�J�a��\���y<>�_/�K%�i�z�g3��S)��U*5-���z'	��Q(�z'	����N�C!��Z�F  ��\'�I��Y�����[�V�B��P�d�i4:=��k5��K%��t-�U*�Z��h�j�J�B���@  0��^��a��\�S����b�d)*��M�s�\'�I$�y<>��o���v�M��y<���?��g3�s9��W+��E�q�|�W+���b��D!(�z����|�o7�M�s9���k��M&3��y<������?��`�t-�����n���r��F��`(4��~�O'�I$����O'�I$��|��w��n�E"1�l�U*5�m��}�?�C�P���I$2�\�g3��F ����F�@�`(4�}>�_��k5��K��I���l���U��z'��d����b���l+������K%�T�e�y��_/�K�R�D�a08��_���u:�^�G�Q�t-+
�R������H"1�l+��E"1�l+�������e2���G#���B  0���O�S��J�B  0�������|��w�].�[��K%�i�z��G#�r��S�T
%)*5�m6�].��m6����k���f�I��Y,6�].7�����N  ���N�C�P$�y<���_�W��j
%)*5���[�V�E"�X�s���G#�r�s�\�����^�A �x�n��A�����C!�h��U��������z�S)*��M�s�\��i4:��O��i���n����h*��M�����O'�I$�y<>?�O'�I$2��N�C�P$2�\�S�T�e�y�~�O'�D!�h*�Z�F�A �x.�[�V�E"�X���i4:�^�G�Q(4���_�W�U�u:=�o7����p�v�����t�V��b$��|���{��O�S�T
%�i��]�w;'	��Q(4�����w�].7�M���|/�K��I$29���k�Z���T��r������X��y<>?�C!��T���Y,�{=�W+
%)�j�e���^�@��P�r������X&������r&3��F�A 08�~��g3��y�~�O��i4:=���{=��k�Z�c1,�{�^�������A�p�v�F�@ �p���m�{=/�K%���E"����C!��T
��I$�y<>?��c��L�Q�t�m�{�^����x����u���_�W+
���d��t-�k����S����b�H"1��[���e��|���{=��k5-���z�������g��l�k5�V�B  08<>�_/�E"�����a����G�Q�����S�T�e�y��_/��e��|�����~�A�p�l+�J!���J!��T
%�i�z�g��l�k��M&3��F���@ �p��[�V�E"1�v�F�A �����c�X�s�\'�I$��|/�E"�����a���N�C��H��Q�t��K%��J�P�d�������i��].7���������a���N��@  08�~��g�Y,6;�N���P�d����b���B�`(��].7���a�x�n��b��D�a�x�n�K%������h�u�����w���W+�J��A 0�|/��A�p��[-��u:=�o�[-+��r�f	���h�u���_/����h�j���Y,6;�g3�s�\��s9��W+
%�i�z�S)�u�}>��o��m6;���c�X&3��F�A�p�l��u�}>��o�[-+�e2����c1��[-�k5���[-+��r�L�c�X�f	��Q(4��~�O'�D����L����\'���R	��Q�������t�m6��n�E"�X&3�L�c���F�A����F��������`(4:�^�������G#�d�i��].��m�{=��w;��s9�w;�N�A�p,���~��c1,6�]�w;��G�Q(����W�U*�Z�����X�����Z���a08<>?�O'��d)�j��E�q�������|��w;���c1�v�c1��[�V�a�x�n��A 08<�?�O'�I$2��N�A�p,�{�^��@��P�d�i�z�N����H���h��z�g�Y�v����i��]�w;�N�@�`(4�}>?���s9�w��n�K�R���A��X�s�\����|��k5���[�V�E��x�n�E"1�l��j��E�q��^�����L���x�n�E"1�l+
%���E"�������X&�Y���m6;����|�W+��E"�X�f�I������e�y�~��@��P��R�D�����F�����B�@�`�h��U*�Z�c1�v�c1��V�a08<������������_/�E"���F�A���L#��R	��Q�t-+�J���`��Z#������P�r���C!��T
%�T
%�T�e2�\����Z�F�A 08��_/�K%���Z����p,6�]�w;'	"1��[�V����P$2�\��i4�}>?�O'�D���X�������f��d��J�B���@ �p�l+�e��|�W���U*�Z���a08<>��o���v��f�����d�T���Y���m6�].7���S)�j��r��S)�u:��O��i��]����~��a0�|���u:�^�C!��T
%��t-+��E��x�n��b$�y�������~���p��V��A�p,6;�N�C!���J�B����D�a0���O�S�T
�R	��x�n�E��x��W�U*5��v�M�s�\'	���h��U�u�}��_/�����T��r���i4���_���u:���g3��F��`�h��U��������z'�D!��T�e���^����X��S��J!(��].7�M�s9��W+��������E��x�n�E"1�l+��r������X&���V��b$��|/�a�x.�[-+�e29�w�].7��f��B���@  ���N��`�t��v���x���k�Z��C!�h��z���c�������X�f	�b��Y,�{�^�C�P��R	��x��W�U���]���}������w��n����������Y�v��f�D�a�x.�[-�k�������Z#�r���i4:=�o�[�V��A 08�~�G#�r��S)�j
��I$29�n�K%�i�z�g3���i4�}>��o7�M�s9.7��h��U�u:�^����@��P$2����c��L�c1��V�a���N�A����F���@  08<>?���q��^�G#��D!�h�j
%���Z��C�P�d�i��]�w�]���}������{=���{�^��c1�l�����n��e2�\�g3�L��h�u�}�?�O'�D�a0�|�o7��f	��Q(4���_/�E���\'�I$29�w;�N�C!������i���n��A�p�l��u�}�������o��m6;���y�~��c1����e�����g�Y�v�M&���V��b��R	�b�H"�X�f�������I���l����j�J��A��X��S�T
�R��B  �x�������n�����l������W�U��z�S��J�B  0�|/�������E�q8���o7�M&3��S)*���f���R	�b$�y�~��g3��S���E"1���K�����I����V�P�����K������d)��U��z�N�C!�h�j�J�a08�����{=/��b��D�P�r&3�f���A���L���x�w;�N�C�P�d�i���n�B�`�h�u��~�C!���J��p�l�k5-�k���f	�q�|�W+
%)���].7���S�T�e�y<������{��O�����M&3�f	���h��U*���f	���h�����j�������J�B�`�h���j���b����A�p�l�k�����i4��~��c1�l�U��z��G#�����`�t�m�{=�o�[��K�R����`�t-+����l�U�u�}>?�C�P�d���Z�F��P������e2���G��h��z���c1�l�U��z��i4�}>?�C!�h���j�J���`�h�u:�^�G�Q��Z�F�A 0��^���q8����w;�������N�C��H"1�v���S)�j
%����M��y�~��g�Y�v�M&3���|�o�����m6;���c1�l�U��z��G��h��z�g����K%)����U*5�V�P�d�i�z�����x����u�}���o7��C�P$�y�~�O�S�T
%�i�z�N�C!���J�����F�@  ���N ��X�s9��W+��E��x.7#��D���D!�t���[����r�L���T�e�y<��?�O'��B �p���K%���Z�Q�t-+�J��H�����J�B�@��P�d��t������[���e�y<>?�O'	"��L����J��A ��\�g����K%�T�e��|�W+
���d�i�����k��M��y�����{=��w�]�w;'��d�i�z�S)*5-��u��~�O�S��J���`(4:�^�@��P$�y�~�����|�o7�M&3�s�\���y�~��g���V�E"1�v�Q(4:�����y<�?�C���D�P$���^�A ����G�Q���M����^��a0���O'��d��J���`�t��v�M&3�L�������c�X�s9��W+��E��x�n��b�H�b��D��p�v��C!(��]�w;�N�C��H"�X�f	��Q(��]����~�O��i�z'	"1,��}�����?�O���t�V�E�q����g�Y�v�Q(4:���g3���C!��T�e�y<����?��g3�L�c1,���~���s9������]���}>�_/��e2��N���������@ �p����v�F��`���J�����H��������x�w�].7����p�l�U*��M&3��S)�����j
%)��z��G#��R�D��H"��L#$2���G#��Y,���~��`(�z�g3�s9���}>�_/�a08<>?��������g3����a�x��{=��w������z��G�Q(��].7���S�����Q(���n���r�f��d�T
%��t���[-�k5�V��b$2�\�g3�L#�����`�h*�����i4:=�o7�F�������A ���N��P�d�i4:���g3�f	��Q(�z��G����J�B ���L��h��U*5�m�{=/�K�R�D!�h������U*�Z�c1�l��u�}���_�W�U*5����m6��n��e��|��k��M���|/���Q�t��v�M�s9.�[��K%��J!(4�}>�_���u�}��?�O'	�q��^�G#�H�b��D�������P��R	�q�����s�\'	��Q��Z��C!(��].7��f�I$2�\���y<���?��g3�L������G��h�j��r��F��`��T�e29.�[����r�L��q8<��_��k5������[-���z�N�C!(�z��i4�}>?�O��i4�}>�_�W�U*5�m6��n��b����A 0�|�o�[�V��H�q8<�?�O'��B �p�v�Q(4:����s�\�S�T
%�i4:��O�S)��U*�Z����\'�I$2�\�g��l�U���].�[-��j��E"�X&��l���z��s����c1�v�c1��[��K%)�u:���g���V��b��D����L�Q(4:��O'����I$29��W�U�u���_/�K%)�u�}���_��k�Z��C!������i�z��G���T
�R	��x��{�^����x.��m�{=�o7�M����^�G#��D��H�q�|���{��O'���R�D�P��Y���m6;��G����J��A�p,6;�g3���|���{�^��c1��V��b$29����u:�^��c1��V���Q(4:=/�a���N�A 0��^���q���O��i�����k���f�I$2�\��i4����o7�M��y<>?��c�X�f�I$��|�W�U���].�������[-+��E��x���������}>�_��k5�m�{�^�C�P�d�T�e�y��_/������V!��Z�F�`(�z�����^����x��W��j�e������s9.����[��K�R	"���F  ��\��i�z��G#�d��J�B��@  0�|�o�[-���U*���f��d�i4�}�?�O'���R	�b���B  ��\�g��l������W��j
�R	������E"1��V��p��[�����Y,��}���_/��p,�{=�o��m��}>��o7����p,6�����u:=����z�g�Y��[-������j�e29�n�K%�i4:=�o�[-�U*5��v��q8<��?������^�C��H"1��V��b��Y����v#��D�a08<�?�C�P$29��{���g�Y���m6��n���Q(�z�S�T
�R	���h���].�[-�k5-���z�N��a0��^�A 0��^�G#�H�b�H��Q����f��B �p,���~��g3���i�z�g3�s�\�g��l��u�}�?�C�P$29��W+�e29���k���f	�b�H�b��R��B �p�l�U*5�m�{=���u:=/��e�y��_�W+�J�B��P$�y��_�W+
������d)��U*5��K%)�j�J�B���@ �p,��}����_/��p���m6;��G#�d)�j�J!�h�u�}�����{��O�S)*5�m6�]���}�?����x�n�E�q8�~��@  �x.�[���e���^�`(�z'	�q���O���t�m�{���g���V�E"������p��V�a�x�w;�g3&3�L��h�u:�^�C�����A�p�v����i4�}�?��a0�|����}>?�C!�h�u��~��g���V���`���M��y��_�W������j�J�P$�y���o7�F���P�d�i�����k5�V�a�x�w��n�K���d�i���n�K%����M&3��F���@���H���\�g3�f�D!��T�����V�E"�X�s���G���T
�R	��x�n�E"�X&�Y,�{����s9�n�E"1�l�U*5�m6;'	�b��R	��Q(�z��G��h��U��z�g3�s�\'����`(���n�K%���Z��q8<>?��c1,6�]���}>�_/���Q(4:=�W+�e�y<>?�C�P$���^�G#�r�L#��D!��T
�R	�q�|�o7����J�B�`��T
��I�r��F���P��Y,6;���c�X�f�D������C�P$2�\�g���V��b�H"1����e2��N�C�P�r��y�~�O'�I$�y�~����D��������H"�X�f�I�r�L�����N��a08<>?�G#�����`���M&3�L#����d)�u:�^�A�p�l��j����Q�t���[����r�f���A��X&�Y,6;'����`�t����m6���W�U�u�}>���w;�g����K�R	��x�w;���c����C!(��].��m6��n���r�L#��Y,6;��s��N�`����E�q8<>��o�������[��K�R	�b�H��Q(4�}����w�]�w;�S�T�e�y�~����x��W+�J�P�r�s9.7#$29.7��q�|��w��n�a�����c��L���T���Y����v�M&����K�R�����P�d)�j�J!��T
%�����Q(4:�^ �������p�l�k5�m6;��G#�H�b�H�b�����R��B�@  �����c���F��`�h��U*�Z�F�A ��\�g�Y,6;�N�C!��Z���a0�|/�K%��J��A ����G�Q�t��K�R�D�a������q���O�S��J!��T��r�f��d�i4�}����?�O'��B�`���M&�Y,6;���c1�l��j��E"�X&3��S)���j��r���C!(4�}����?�O��������i�z�g�Y,�{��O���t�������m���~�O���������t�m��}��_/���r��y<����o�[-+���������b��R���A��X&���V���`�t�V��A �x�w���W+��E���\�S)�j�����h�u:�^���q��^ �p��V�E�q�|���{��O'�I�r���C!(4��~���s9.��m��}>���w;�N����X������g��l��u:=��k5���e2�\�S)�u:���g3�f	�b�r�s9�����_����z�g��l���U�u�}���o7�F������A�p��[�V���`(4:=��w;�N��a��\'�D�a0�|�W���U�u:=��w;'	�b��D�P$��|���{�^�G��h���j
�R�D�a����G#���B���H�b�r&3�f�I�r��F�A�p��V�E"���F�`�h*����S��J�B  �x.��m6;�g3�f�����d)�j
���d)���j��r��F���@�`��T
��I��Y,�{��O���t�V�a0�|�o��m�{=��w;�g�������Y,�{=����}>?�C!��T�e2�\���y<�������{=�o7����p,����_���u�}>��o7��f�I�r��S��J��A ��\���y<>��o7��f�I��Y,�{=/�K%�i4�}>?���s�\���y<>?�O�S)*5���[-��j��r�L�Q�t���[-�k5�m�{�^�G#��R�D!������Q��Z�F�A��X�f	"����C�P��R	��������Q(4:=/��e�����g��l�k����S����b�H�b�r��F��P$2�\��s�\'�I$2��N��a08<>�_/���r�L���x.��m�{��O�S)�j�e29�w�]�w;��G#�d�i4:=��w;��������s9���k5��K��I�r�f��d�T
%����M�s9.7��C�P��Y�v�F�A 0�|�o��m6;�g�Y���m�{=�����~���s9�w;�g3�L��q��^�G#$�����g3�L#$���^���p���m��}���o��m�{=/��A�p�v�c1,��}>?�������G��h�u���_/�a������q8���o7��f	��x��W�U��z��G#�r����a0�|/�K�R��B���H�b�H�b$29�����z��G���������T
%��t�V����h���������j
��������I�r���|�o7���������S�T
%)��U*�Z�F��`(�z������O'�I$29.�[-���z�N�C!�h�j�J!���J!�h�j�J!���M&3���i4:�����y��_�W+�������e��|�W��j
%�i�z�N��a0��^��c�X�f���A 0��^��c�X�f�D��p��[-+���b��D�a��\'	�b�����`(4:=�o�[���e2�����q8��_/��e�y��_�W���U*5�m���~���q��^�G#��D!����f��d)*5-��u:��O�S)���]��{��O�S��J��A �x����u��~�C!(����W�U��z�S��J��A 08�~�O�S����b�d)����U*5�m6;�g3�f���R��B�@�`������Q(4�����w��n�K%���Z�Q���M���|�o7���S)���]�w;����q��^�A 08����������w���W+�J�P�d���E"���F�`����E��x.7���S)�u�}����w�].�[-�k��M�s9������o�[-+���b$2��N�A 08<��?����y�~�O'����`��T�e����O��i�z'	���\'����I$2����c�X&��l�U*5�m6;�����^�C!�h*5����r�f	"�X�f��d)��z�g�Y,6�]�w;�S��J������D!�t�m�{=������_/��p���m6��n�K��I�r�����p�v�c1�v��f��d������S)���]���}>��o7�������F�`��T
%���E��x.���v#�d)���j�e��|��k��M&�Y���m6�]���}�?������N�A�p�l�k5-��j�e��|���{�^�G���T�e2�\�g3���C!�h*�Z��C!�h�j�J�a0�|���u:=���u�}����?����x.��m6�]����~���s���G#�H�b$29.7���a����G#�r&�Y�v�c1��V�B�`(�z������f	��Q�t�m6�].7�M&3�L�Q��Z����J��p����e�y<���o7�F�A��X��S��J�B����@  �x�n�K%��t-��j������T
%��J��p�v�M&3�f	��x.�[��K�R����`�������h��U��z��G�Q(�z���c��L�c1,�{�^  ���N�C!�t���[�V����h*5-�k5-���U*���f	�b���B��@ ����F�A��X�f���A���L���T
%�i�z'	"1�l���z�N���p,��}���o��m��}>?�C�P�d)�u:=/��A 08��_��k��M&�Y,6;����Z#�d�i4:��O��i4:���g3&3�L�c�X��S�T
�R	"1����v�c1��V��A 0�|�����~��g3��F���P��Y���m6;����q8���o���v��C!�h������U���]�w;����q��^�������A��X���i4��~�G#��D�a�x.7��h�j����Q(4:=������_/��e29.��m�{=�o������v��f�D���D���D!���M&��l����]�w;��G#��D�a�����c��L�Q(��]�w��n��e��|/���`��T
%��J�a��\��i��].�[���e�y��_�W�U���].7���a0��^��a���N�����D���X����t-+���b���l���U*�Z�F���P$�y���o�[-��u:=/!�h*�Z#���I�r�s9��W����j
%�T���Y,����_/���r�L���T�e���^�G���T
%�T��r��F���@  08�~��`(���n�a08<>?��g3&3�f��d��t�V�B  0������y<�?���s9�n��b�H��Q(��].�[�V�a�x.�[���e2�\�S)��U��z��i4:=���u:��O�S)�j�J�B��P���I$29.�[�����Y,�{�����y<���o7���T��r�����p�l+�J�a�x�n���r��F���P�r�f�I$��|/�K%�i���n��b$�y<>?�G�Q�����S���E"1,6���W�U*5-��u�}�����_/�B�`�h*5���[-�U���].7�Q(4��~�O��i��].�[�����Y,6;'�I��Y�v�M&3�f	"�X��y<>�_�W+
���d��J�������B ���L��h*5��K%)*5-���z�N��@�`��T�e�y�~���s9���k�Z����\'��d�i4���_/�������K��I$2�\��s�\��i������u�}��?���s���G�Q��Z�F�`(��]��{=�o�[-�U�u�����w;'�D��H�����G#�d�T�e�y��_/�a0���O��i4:=����}>�_/��b���B�@�`�t-+�����h�u:�^�G#������I��Y�v�M&3�L�Q(4�}�����o��m��������}����_/�K�R	�b�d�i4:���g���V�E"1���m�{�^�@��P$29����~�G#�H�����G#�H�b��Y�v��C!(4�}>?��g3&3�L#�r��S)*�Z�F�A 08�~�A ����G#���I�r�����p��V���`(��������].�[������l��u:����s9.7�F  ����G#�d�i4:=�o�[-��u:=/�E��x.7����p,�{=��w;�N����X���i4��~���q�|�o7�M&�Y,6;��G#��D����L��h��U*5��v��h�u:=/��p��[�V�E"1��V�E�q��^��a08<>?�O������f�����P�r�L���x��W�U��z'��d��t������l+
%��t-���z�N  08<>�_�W+��r��y<>����{�^���@�`���M�s���G�Q(�z���c���F�����@�`�t-��u:�^��c1,6����k�Z��C!���M&3���C!��T
��I����V!(��]��{������|/��e�y<>?��@���H�b$29�n�K��I$�y<>�_�W���U�u�}>?�O�S�T
%�i4:=�o�[-�k��M&3�L#$�y<>�_�W+��r���|/��A �x������].7��h*�Z#�H���\�g����K%�i��]�w;'���R���A����F�A��X�f��d��J����L�Q��Z�c1��V����h��U����n����h�j�e�y<��_/!�h�j�e��|�W����j�J�P�r�L#�����`(4:�^���p�l�k����S)�j�J�B�@��P�d����M��y<��?�G��h��U����n���r���C!(4:=�o�[-���������z'	���h�j
�R��B �����C�P��R�����P�����R	�b�����`��T��r�����p�����r����a08��_/��e29�w;�g��l�U*5���[���e2��N�@���H��Q(�z�����x��W��j
%�T
%�i4��~��g�Y�v���S)*5��v�M&3�f�I����V�a08��_/��e�y��_/�����l��j��E��x���k�Z�c1,6;�����M��y<>?�C���D�a�x�n�B  �x�n�E�q��^��c��L#��D!���J�B��P�����R	��x��{=�o��m6�].��m6;�N�@ �p�l������j��E�q�|�o7�M�s9���}�?�O��i4:��O����Z�Q��Z#��R	�b����A�p�����r&3��y��_/�K��I�r��F��`�h�j�e2�\��s9�n�E�q8��_/�B������A�p���m6�]�����_/��e�y���o7��C�P$29���}���?�O'��d��t-��u:=�o7�Q(4:�^  ��\'�I�r���C!(�z�����x�w����k�Z�F�@ �p,�{=/���`�t�m6;���c1�����r�����p�v�M&3��F���P��R	���\��i4:=����}>?��g3&���V!�h*5��K�R�D��p���m�{��O'	���\'	�b��Y,�{���g�Y��[-�U�u��~�������O'�I$29�w�].7#��R	"��L#�H��Q(�z�g3����a�x��{=�o��m�{��O���t���[-�k5-�U���].7�F����H���h�j��E������c1���m6;�N�`���J�B  0���O'��d�i�z���c1�l��u�}��_/!(4�}>?�O'�I�r���C��H��x��W�U*�Z��q8<>�_/�K�R�D!�h�j�e���^�G�Q(4�}>?�O���t��v�F�A�p�v���a08<������_�W+�J�P����d�T
���d�i�z�N�`(4��~�C!(�������z��G#��R	"1,�{�^��c1,���~�O��i��]�w;'	�b$��|�����~�G#�H�b$��|�W+���Y������m6;�N�����L�c�X�s9�n��e29��W+��E�q�|/�B�@ �p��V�E��x��W�U*5��v��h��z���t�m6;�N���@  ���N���p�l���U*5-��j��r�L�Q��Z�F�A �x�n�������E�q8��_/�E"�X�s9.��m�{�^��c�X�s��N�A ��\�g3&�Y�v�F��`�h���]�w�].�[-+
��I$29.����[-��j�J����P���I$�y<������w�].7�M&3&�Y,6����k���f�D!��T
�R	���h�u�}�?��g�Y,6;'���A 08�~�C!���J!�h��z'	��Q(��].7�M�s��N�C��H�b���I$��|�W+�J��A�p�v��f��d�i4:��O'�I�r���C�P$��|/��e�y�~��g�Y,6;�S)���j�J�a0�|/�K%�i���n���X��S����b����d)*�����i�z�N����X�f�I�r�L�c�X�s9�n�K%�i4�}�����?���s9�n�K%)�j���b�H��Q�t�V�a08<>���w���W�U���]�w���W�U��z��G�Q��Z�Q����f	��Q�t�V�E"���F����@�`�h�j
%)*��M�s9�w��n�K%�i4��~������^�G����J��H"1,��}���������}���_��k5��v����p�v��f��d�i4��������~��g���V��b�H����T�����������V��A������a������q8�~�O'���R�D!��T
%�i4�}�?���s9�w�]��{=�o�[-�k��M���|/��e��|/���Q(�z�N�A 08<>?��c1���K%�i�z�S)�j������T���Y�v�M����^�G�Q(�z����Z��C��H��Q������i�z�N�@  �x�n��b��R	�b�r����a��\'�I$29��{���g����K�R�D��p��V�E�q�|�W�U���]��{�^�G#��D!(���n�K�R��B �����������C!���J��A �x�w;�S���E�q��^�G���T
%������h�u��~��c1,6;�N��P�r��S���E"1������Y���m6�]���}�?�O'��B �p�l+�J��A��X�f����`������������Q(�z��G#���I�r�L�c��L�Q�t�m6;����|/�B�@  �x���k�Z����\���y��_���u�}�?�O'�����d�i4�}�?�O��i4�}>����{�^���q8�~�O��������i�z��s��N�A ���N�C!��T
�R	��x��W+�J!�h*5-��������u:�^��c�X���i��].�[-�k5-�k5��K���d����b�r&�Y,��}��_��k���f��d���E"1�l�k5�V�P�r��S)�j��E�q����g���V�a�x�n�E�q�|���u:=��k�Z�F������@��P�d)�j���Y,�{�^���P$29.7���S)��U�u:=��w�].7������G��h*5-�k�Z��h�j�J�a�x.�[�V��A���L�Q��Z�F�A �x���k5����m6�].7���S�T�e�y<�?�O'��d�i4�}�?���q8��_/��b��R	"1�v�M&�Y,6;'�D!(��]�w;�g������r�f�D��H"1�l+�e2�\�g3����a��\���t�V��A�p,6;����q8<>�_�W��j����Q��Z��q��^�G#�r���|���u:=����}>?����y<>��o�[-�U*�Z��q8�����{=/�E"���F���P�����K%���E"1,6;����q��^�C!(4�}>?�O�S)*��M&3&�Y��[-�k���f	�b$29��W+�J!�t-�U*5��v�����t-�k5��K���d)��U�u��~��P$�y<������w��n�K�R�D!�h*5�m6�].7��q����g���V�a�x.�[������l�U�u��~�O'������R	����T�e2���G#�d�T
��I$�y<>�_/���r&�Y��[��K�R	"1�l+�J�P��R	�b�H��x.�[-�������k5�m�{��O'	"1,��}>�_���u�}>����{=��w��n��e���^�G�Q(4:�^�G#��R	�b�H�q8<>�_/��b�d��t���[-�k�Z�c1,���~�C�P���I$�y<��������_������n�E"��L�c1�v����i4:=��w;��G#����d�T
�R�D�P$29�n��b�H"������p���m��}�?�O�S)��U���].7�M��y�����{�^����x��W+
�R	��Q(4:��O'	"�X&3�L�Q����f���R�D�a�x��W�U*�Z#�d�T
%��J����P�r�s9��{�^��c1,6;�N�����L����\���y�~��a08������}�?�C!�h�����W+�J�a�x�n�K��I�r���i4�}�?�O'����I�r�s��N���P�d�T
��I$�y�~�O�S)���].��m6���W+
%)�u:�^����X���i4:=�o�����m�{�����y<>���w;����Z#$�y��_/��e2���G�Q�t�m6����k��M&����K���d�i�z�N���p�����r&3���C�������P��R���A�p,���~����y<����w;���c1,6;�g3����a08<��?��c�X�f���R	���h�u:=��k�Z�c�X�f�I�r�����p,��}�������?���s�\'��B����D���X�f	����N�@�`�h�j�e29��{=�W+
���d�����Q(4��~��g��l��j�J��A 0�����s9���k5���e29�n�B ��X�f���A�p,6;�N  08�~��P$��|�W+�J!�h�u�}�?�O��i4���_�����]���}>�_����z��G�����E�q�|���u�}>���w��n����h����U*5-�U*��M&3&�Y�v��f��d��t-�k�Z�Q(4:=�W�U�u:=�o7��f	�b�d��J!�h�u:��O�S)�j���Y�v��h��U*5�m�{�^��c�X��������S���E"1����e29���k5��K%���E"�X�s�\'	�b��R	���\�S��J�B�`�t��v�M&��l�k5��K%��J���`�t-���U���].7����i�z��G���T��r���|/��e�y<>�_�W�U*5�����Y��[�V�����T
���d�i�z������\���y<>?�G������b$29�n�E����N�C!�h�j�e29��W+�e2�\'�I�r�f�I$��|��k5�m�{�^�C!��Z����J����L�c�X�f	�b�H��Q(4���_/����Y,���~�O'�D���D��p��V�a08<>�_/����B�@ �p�l��������j
��I��Y,�{=/���`��T
�R����`���J�B  ��\�S�T�e�y���o��m�{�^��c1,�{���g3��F��`���J���`(��]��{=/!��T
�R�D!(�z�N�C��H���\�g���V�E"1��[���e29��W+��E��x��{=�o����[-����j
%��J�a0�|�o����[��K��I������e�y��_�W+�J!��T��r����t-+�J�B��P�d��J���D!�h*�Z�F�@  �x�w;�g3��S���E"1,���~�O�����M�s9���k5�V�����T
��I�r�f�I$2�\�g�Y,�{�^�C�P�r��S�����Q�t�m6��n�E���\'�I$2�\��s���G�Q(4:��O'�I���l�k5-��j��E"1,�{=�o����[����r&�Y,�{=�o��m��}��_��k5�m�����o7�c1���m�{=�o7�F�A 0��^�A 08<>?��g3�f��d�i�z�g3���C�P$����O�S)�u�}>�_/�E"�X&3�f�I�r&3�f	����T
%)�j
%�i�z�����x��W�U*�Z�c�����a�x��W+����l��j�����h��z'��d�T���Y,�{=/�K��I$��|��k�Z���x�w�]���}����������o�[-�U*����S�T
%��t����m6���W�U�u:���g3��y�~�G#����d�i4��~��g��l�U���].7���a��\'���A 0��^�G���T
%��J!�t-��u�}��?�G#��D��������p����������e��|�o7�c1,6�]���}>?���s9.7�����t�m6;'�I�r��S)�u�}>?��g3�L�Q�t-���z�N��a0��^����x��W+�J�B�@ ��X��S���E"���F��@�`�h�u�}���o7���S�T
��I��Y,�{=�o7�M&3�s9��{=/���Q������i�z�S�T
%�i4:�^��c1��V��p��V�E����N�A ��\�����M&3&�Y,6�].7�F�`��Z�c�X�f��d���Z��q�|��w���W+����Q��Z�F��`(4���_/�K�R�D�����F�A 08<���_�W��j��E�q�����s9�n��b��D�P�����K%��J�P���I$��|/�K���d���Z#�d��J��A 0�|��w�].�[�V�E"���F �p�l+�J�P�d)�u��~��c1���m6��n�K%)��U���]��{=/�����H�b���������I$��|����}��_�W�U*�Z��C�P����d)�j�e29�n�K%)*5�m6���W+�J!(4:�^��c1,6��n!���J�B���@���H��Q�t�m��}���?��g3�L#$29�n�K%�i�z��s9��{���g�Y�v�F���@ �p,�{�^��a�x�n�P���I�r&�Y,6�].�����m��}>?�O'	"1,6;���y<>?�O�S��J������`�h*5�m6��n�K%�i��].7���S)���].7#�d�T�e2�\'	��Q�t��K�R�D!�h�u:=�W�U����n�����������F�`�h*5�m�{�^�G����J!�t�����v�M&�Y�v�M&�Y��[��K���d)����U*5�m��}>?�G#$29�n��b$2�\�S�T
�R��B��P��R�D���D�������a0�|������n���r�L��q�|�o7��f��B ��X�f�I$��|/�E�����G��h�j�e2�\����Z�c�X��S)*�Z#������I$2��N���p,�{���g3�s9���}���o7�c�X���i�z�N���p,�{=�o7�M&3�L#���l�U*�Z�c��L#����V�E"�X��y<�?��c�X�s9��{�^��c1,6����k5�m6;'���R	�q8<>?��c�X��y<>�_/�E�q�|�o7��f�D!����E����N�C!(��].7�M�s�\�g��l��u:�^�G�Q���������M&3���C�P�d�T
%�i4:�^�G��h��z�g��������l+
%)�j����l���U��z�����^�����D���D!��T
���d�i4:=/�E"�X���i�����k5��K%��t���[-����]�w;���c1�v��f�I$29���}>�������_�W��j
%�i��].7�F��@�`(�z��G#���B �p��V�E�q8�~�G#��R��B��@��P��R	�b$�y�~�����\�S)��U*�Z��C!(4:�^��a�x�n�����l+�J�B�@���H�����J�a�x.7������L��h���].7����i�z�����x.���v�F��`�t��K�R	"1,6;�N  0��^���p,���~���s9����u:=/!(4:=�o�[�V�B�@��P�d�T
�R	��Q�t���[�V���Q(4�}��������~�������@���H"1,�{�^��c�X�f�I�r�s9�w;�S)�j�J�B  0�|�o��m�����o��m6���W+�����h*��M&�Y�v��C�P�d�i4��~��g3����t��v��h*5-+�J���X�f	�q8<>?�G#�H"��L�c1��[-�k5-�k�Z�F�`��T�e29����u�������}�����w����k��M&3�s��N���������P����������V�B��@�`�h�j��r&�����e29��W�U�u:=��k�Z�F�A 0���O�S�T�e29����u���_�W+��E"1�l��j����Q(�z��G#�d����M�s���G�Q(4:=��w;��s�����q���O��i4:�^��c1�l���z���c1��[��K%�i�z����Z���a08<���o7�M&3�L����\�g���V�E"1,6��n���`�t�m�{�^���p,��}�?��c1�v�����N�@  08<�����o�[�V����L�c��L�c���F�`��Z��h��U���].7�F�`��T����l����j���b����A�p,6;���c��L#$29�n�B�@  08���o7��C��H�b��D!(4:=�o7�M�s9�n�K�R������H�b�������������H�b��Y��[-�U*5-�k��M&3�L�c1�l��u:=��k��M&3�L��q����g3���C��H"�X���i4:�^�G���T
�R�D!�h���j��E����N �p�v�Q��Z���x�n�K%)����������U*�Z�F�A�p�v��f	������c1���K���d)�j��r�f�D!�t��v��C����B�@ ��X���i����W����j�e2�\�g3��F�@�`��Z�Q(4:�����y<�?�C�P�r�L#�H�b�H���h*5-���z���y<>�_/�E���\��s��N�`(��]��{����s9���k�Z�����X&�Y���m6;�N���p�l�k�Z�Q(4:=�o��m6��n���������Q����f	"1�l�U*�Z������L�c�X�f	���h�u:���g��l�k5��v�F�A�p�l�U��z���c1�v�M�s��N�`(4��~���s9��W��j
��I$�y����w�].7��f��d���E�q�|/�K%��J�B ���L�Q(4���_/���Q��Z�Q(���n�K�R�D�P�d����M��y�~�C��H�b�d)�j�J���`(4:=��w�]�w;�N�C!�h*��M&�Y,�{��O�S)��U*��M&3��S)����U���].7�M&3���C��H�b����A 08<>���w�]�w;'�D!����E�q�|�o7�M&���V�E"1�l��u:=/��b�H��x�n��e2��N  08<>?�O������f��d�T
������d)�u:�^��c1,�{���g�Y,6���W+��r�L�Q�t�m6;�N�`�t���[�V�a08�~�C��H���h�u:=/�K��I$29�n��e�y<>�_/��b���l��u:=�o7�F�@  �x��{�^�����\�g3�L���x.��m�{=/!(�z���c�X�f	�q8<>�_/�E�q8<>��o7�M&���V�a�x�n�K%��t���[�V��b�r��S��J�B  0���O�S)�j�J�B��@��P$�������y<��_�W�U�u�}�������}��_/���D�P���l���U*�Z�F�@�`�����b�����`��Z�F���P��R	"�X�f��d��t-+�J!(4:�^��@  �x��W+�J�B�����@  0�|/���r&��l+��E�q��^�C!�h�j
%)�u��~�O'	�q��^�C�P�d�i�z'�I$29����~���p�l�k5-�U*5-�k5�m6;�N��P�������d�i����W����j
�R	"1��[-��u:��O'��B��P�d)��U�u:=/�K�R	��x��{=��w;�N�@  ��\�g3��S�T�e�y<>�_/��b$2�\��s��N��a�x��W+
%�T
%��t�m6;����q�|����z��s��N�@��P�d)����n���r�L�c�X�f	�q����������g3&3&�Y��[�V�E�q�|��k5�m��}��?���s9���k5-�������U*5-�U�u:=�W+���b$29��W�U�u:�^�G#$2��N���@�`���J�B�����B�@�`�h*���f�I��Y,6�]���}>?�O��i���n������V�E"1��V�E"1��V��b��D����L��h�u:�^�C��H�q8<����_����z'���A ��\�S�T
%���Z�F���@ �p��V���Q�t-�U*5�m��}>���w;��G#�H"1,6;�N ���L�c�X�s9�w���W+��E�q8�~�O�S)����n�a��\�S)���j�J!��T�e�y<>�_/�a0��^�G��h�u:���g��l��������u��~���s���G����J��A 08<���?�����|��w;��G�Q�t-�U*5-�k�Z�F����H�b��R�D�a0��^�G�Q(�z��G�Q��Z�c�X�f�I$�y���o7��C��H��Q(4:=��k�Z�F�����D�a0���O'�D�a08<��_/�E��x��W�U��z'�I$29�n�E"�X&�Y�v�F  08�~�O��i���n��e2���G�Q�t��v��q8�~��c��L�c1,�{=/�E"�X��y���o7���S��J�a�x��W+
%����M���|/�K�R	�b���l+���Y������m6�]�w�].��m��}��_���u:��O�S)���]�w�]�w;��G#���B���H�b�r�f�����d��t-��j�e���^��c��L#���B  �x��W��j�J�a0���O�S)�u:����s9�w;�N�C!��T
%)���j�J!���M�s9�w�]��{=���{=���{=/�E��x�n�K%��t��v��f�����d)�j�e2���G���T��r�f�I$2�����q��^�C������`(��]�w;�N��`�t�m��}>��o��m�{=����z�N��@�`��T�����V�E"��L#�d)��U�u�}���_/!����f�I$����O'�I$2�����q��^ ������a0����g����K����R	��Q(4:=�o7�M&�Y,�{=/��e2�����q8<>?�O'�D��p�v�M&���V�B�@��P��R	�b�d�T����l��u����o�[-��j�J���`(�z�g�Y���m6���W���U*5���[����r�s��N��a���N�C�P�d)�j
��I$�y<�������~��c1��V��b�d���Z�Q�������t�V���Q(�z'�I$2��N�@  �x.������v��f�I��������Y�v���a��\'�D���X��S)���j�J�B�@���H���h��U����n��e2�\�g��l+���Y,6;�N�@���H�b�����R�D���X�f�I��Y��[��K%�i�z�g3&��l��u���_/�E"1��V�E�q8<>��o7�c1�l�U��z�g3&3�L�c���F��@��P$��|����}>?�G�Q��Z�F�@ �p,6����k�Z#��R	��Q�t-+�J!(4:=�W�U�u:���g3��y<>��o�[�V�a0���O��i�z'�����d�i�z�N�������C�P�d��t-�k5-+�J�B  �x��W�U*�Z���a08�~�`�h����U*��M&��l�����n�B���H"1���K%�i4�����w;�����M&�����e29��{����s��N���p�v��h�u:��O�S)���j�J�a0��^��c1���K���d)��z�N���p�v�M�s����c1��[���e2�\'	��Q(��].7�����X����t�V!(��]��{=��k��M&3�L���x.�[��������K%��t�V���Q(4:=/�K�����I$2��N���H"1�v�F�`�h�u��~�G�Q�t�����v�M&3���i4:=��w��n�a���N�C����B��@����D�a�x��W+
%)���j��r����a����G#�d����M&3��F���P�d�i�z�g3�s�\�g���V�B�@�`�h�j�J��A ��\�g3&3�L��q���O'��d�i4:��O'��d�T���Y,6�]��{��O'�I�r���|/�B��@���H��x�n��e2���G�Q�t�m6�]��{=�o7�Q(4:=/�B  ������q8��_/�a�x.��m���~���s��N�C��H�q8�~��g��l�k5�����v����J�P$2���G#$��|�o�[�V����h�u�}��_��k5��K%�i4�}>?��c�X&3���C!�h*5��K%���E"�X�f������R	�b$���^��a08�~��c1,���~�G#���B  0�|�W+���Y��[-���U*�Z�Q(�z��i4:=��w;�g3����a0�|��w;�����x����u:�^��@�`(4:�^�C!����E"1��V�B�@ �p�l+
%��t�������V��b$29��{��O'�I��Y��[-�k�Z�F�@�`�h*��M&����K�R�D!����E���\�S)���j��E"1�v��f�D���X�f�I�r���C���D������`��T��r�L#�H"1�l���U��z'	����T
%�i�z'�I�r&3�L��q�|��w��n����P�d)��U�u:�^��c��L����\��s��N�@�`���J��p�v���S��J�B �p�l+��E"�X�f�D��p�l�U�u:��O��i�z���c1���K�R	���h��U*�Z�F������B ��X�s9.7��f�D�P����V���Q�t��v�M�s9�w����k���f�D�a0�|�W��j�J���X�s���G�Q�t�V�E"1�v����i4��~����H�b�����K%���Z�Q(����W����j��r�f�I�r����t��K%�i�z�N�@  �x�w�]���}��_�W+
���d�i4:�����y��_��k5��v�M�s9�w���W+���b�d)�u:=�W�U*��M��y����w;�S)��z��G#���B �p���K��I�r���C!��T�e2�����q8<������}��_�W+
��I�r�s�\�g3��S�T�e2�\���y<���_�����].7�M����������^�G#�H"�X�s9�n�a0�|�W+�J��A ��\�g3�f�D��p��V�E����N�A �x�n�E"�X�f���R�D���D��p�l�U*5��K���d���Z�Q�t�m6���W���U*�����i���n��e2��N��a���N��a�x��{=�o7�M�s�\��s9.7�M&3�L#$�y<�?�����|��w�]��{�^�G�Q���M��y<�?����X�f�D�����F���P�d)���������]��{=/�a08�~�O���t�V������������J�P�d��t�m��}>��o����[�V�E"1��[���e�y��_/�B��@��P�r����t�m�{=/��b$�y���o��m6��n���r���C��H�b��R��B�@  ��\��s��N�C!�t�V�B�`�h�j�e�y�~��a�x��{=�W�U���]�w;�S�T
��I�r����t�m��}>?�C!�h��U*�Z�F�A 08<�?��c1�v�M���|/��b�����R	"�X�f�D�P�d��t-������j����Q(4:=/�K�R	����T
%���E��x�w;��i4:=�o�[-���z'	���h*�Z��C�P��R��B�`���J�B ��X��S)���j�J��A ����G�Q���M��y<���?��a08<>���w�].��m6;�S)�j
���d)��z��G#$���^���P$�y��_�W����j�����V��b��R	��Q����f	"�X�f	��Q(4�}�?��g����K%�T
%�T
�R	"����C!��Z�F�@  �x�����z�g3�L#�r�s9�n���Q��Z�c���F���P�d�i�z����|��k�Z�c�X��S)���j��E"��L#��D���X�f�I��Y,�{����s��N��P$�y�~�����D!�h�j
��I$�y�~��g3�L�Q(4:����������s9��W�U*�Z���a��\�S�T
���d)���j��E�q����g3��S�T
�R	���\���t���e��|�o�[�V���Q(4��~�C!�h�j
�R	��Q����f�D�a08�~�O'�D�P��Y,6;�g3�������L#����A�p��[-+���Y,�{=/�K%�T��r����a08�~�O'���A �x�n�K%�i4��~�O'	��Q����f	�b�r���C�P�d�T
%�i�z'����I$2���G��h�������j���b��D���X�s9�n��b��R����`��T���Y�v�M&��l��u:=/��A 0���O'��d���Z���a0�|/!�h���j�J�B��@  �x��W+���b�H�b�H���h��U*�Z���������a0�|�����].�[����r���i�z��s9.7�M�s�\���y�~��g3�f�D!��T
��I�r�f��B�������@�`�h�j
%����b�d�T
%�T��r�L����\���y�~�A ��\'��d���Z���x��W+
%�T���Y,6���W+�e2���G���T���Y����v�M&��l�k��M&��l��u�}>�������_/�K�R	��x.�����m6;�g�Y,���~�@ �����C!��T��r�f��B �p�l�U�u�}���?���q��^�@�`�h���j
%�T�e����O���t-��j��r�f���A������a0�|���{����s9�n�������K�R	"���������F�A�p,����_��k�Z�c1,6�].7�F �p���K%)�j�J�P$29��W+�J��A 08<�?���@ �p��V��b���B  0����g��l��j�e��|���u�}����_/�K%�T�e29.��m6�].��m6�]�����_��k��M&��l��u�}�������?�O��i4�}>�_�W��j�J����L#$��|���u:=/��������b�H�q8<�?�O��i�z�N�@�����B�`�h*5�m���~����X��S)����U*5�m�{�^�C��H����N�C!(4:�^�G#��Y,�{=��w;�N�@  08<>�_�W�U*�Z#��D�P$�����g��l�k5��K��I$��|��w��n�K���d�T�e�y���o7�M��y<��_/�K���d)�j�J�B�`�t��v�c1,6;��G�Q��Z������������L���x��{=�W���U��z'�I�r����t�m�{=�W+����Q(��].��m�{���g�������Y,���~�@���H���h�j�J��A��X���i4�}�?��c���F�`(4:�^�G�Q(4:�^�G�Q(�z�N�C��H"����C!���J!�t���������e��|�W+�e2�\�����^���q��^�A �x.7#�H�b�d��J������������D��p�v�c1�l�U���]���}�?�O�S�T��r�s9���}�?�G#���I�r�L���x���k��M�s�\'����I��Y,���~�O�S)�u:�^�C!�t�m�{=/���r��S)����U���]�w������������z����q8�~��g��l�k��M&3&��l+�J���D!��T
%)*�Z�F�A �x�w�]�w;�S)*5-+���������b���I$���������^��c�X&3��S�T��r�L�c���F  �x���k��M�s�\�g��l�U����n!����E��x��{=�W�U��z��G#��D!(���n��e2��N�C!(4�����w�]�w;�N�����@���H�b�H���h���]�w��n��e�y<�?��c�X&�Y���m6;�N�C�P��R	�q8�~�O'���R�D������C�P�r��F�A�p�l+�J���`���M��y<>?���s9��W�U��z�g3�s9���}�����{��O'	��x��W�U*�Z#�r��S)�j�e��|��w;�g3�L��q8<���o�[�V�E"1�v�M�s�\'	��Q(4��~�O'�I���l���U*�Z�F�@���H������E"1�l���z��G#��D�a��\���t-+
�R	"1�v�c�������X��y��_/���r�L��h*�Z�F  �x�w��n��e29.7�M&�Y,6�].��m6���W+���Y�v��q��^�G#$2���G���T������K%�T�e���^�@�`(�z�N���p�v��f��d)*�Z��h�u�}��_/�K�R	���\'��B��@�`�����b�H"�X�f�I��Y�v��q�|���u��~������N��`�h��U��z��G�Q(4:�^��c1��V���Q��Z��h*�Z�����X�f�I���l�U*����S)*�Z�F  ��������\�g3�L#���B ��X���i4�}>�_�W���U*��M�s9��{�^�G�Q(�z�N�A 08<�?�O'��d�i���n��b�H�b��Y��[��K����R	"1��V�a0�|��w;'���R�D��H�b����A�p�v���a���N�`������i���n�E�q���O�S)�j�J�B��@��P��R�D����B��@ ��X��S�T��r�L��h*5�m6;����Z��C����B��@  08���o��m6�]��������{�^�@�`�h�u:��O'�I�r&�Y,�{=�o7��f��d��t���e���^��@ ��X����^��c�X&3���i4�}>?�G�Q���M&3���C��H����T��r���C�P�������d���Z#����A ��\�g���V���`(4:��O'	��Q��Z��C�P���l+�J�a��\'��d���Z�F����H�b�H��Q��Z�c1��V����P��R	�b�H��Q�t��v�F�A�p,�{�^�G�Q���M&3���C!��T��r��S)�j��r���i�z�g�Y,6;�S)�u�}��_/���`(��].7�F�A ��\�S�T�e���^��c�����a�x.�[-����j���Y,6;���c1�v�M��y�~�O�S)�������j��r��y��_����z�N����X�f��d)�j
%�i4:=�W����j�J�������P�d��J��A 08�~��g��l+�J!(�z�S�T
%�i4:=/�K%�i��].7�F�A 0����g3��F�A 0��^�G��h*5-�k������t�V�B�`�t�m��}��_�W+
����������R	"1�l+��E�q8�~���P���l�k5���e29���}>��o7�F�@ �p�v��f����I$29�n��e2�\��s9�n��e2�\'���R��B���@ ��X��S)����U�u:�^����x���}�?�C!�h�u:�^���q8�~��c���F�A�p��V�E"�X�f	��x�w��n�K�R	"��L�c1�l���U*5��K�R�D�a��\��i4:=���u:���g��l�U*5��K%)*���f��d���E�q���O�����M&3��y�����{=/��b$29��{=/�E"1��V���Q�����S)*5��K%��J!�h�j�J!�h*�Z��C�P$29�n�E����N����X&��l+���Y�v�Q(���n�E"1���K��I$�y<�?�O'��d�i4�}>?�G���T
%�T
%���Z��q����g3���C!(4:=��w�].7��f	�q8<�?��c�X�f��d���Z����p��V!(��].7����p���m6;'	��Q�t���[-���z�N�����@�`�t-���U*5�m6;�N�C�P�d���Z#$������s����c�������X&3�s9���k�Z�F�@���H"����C��H��Q(4:�^��a��\�g3�f�������D��p���K%)�j�J�����F�A��X�f�I$29.7��f�I$��|�o7��f��B�����@�`��T�e29�n�E"��L�����N�@  ��\'�D�P��R	�b�H"1,���~��c1,6;�g3�L�Q(����W+
��I$�y��_/�B �p�����r��F�A 0�|/��e2�\�S)��U��z��s9�n�E"1��V�B�@ ���L#�H�b����d�i��]�w;�g�����e��|��w;�g3&3��S)*�Z�F��`(4:�^�G#�H"���F��`�h��z�N��@�`��Z�������F��`�h��z����|/�E��x�������w;���c��L�c�X����t��K%��t�m�{=�o��m6�]�w��n�P�r��F���@ ���L���T��r���C��H�b�H���h��U*�Z#�r��F�@  ��\���t�V�E������c��L�������Q(4:=��w��n�E����N����X�������f��d���Z�F�A �x�n�K��I��Y�v�M����^�G���T
�R���A��X�f�D����B�@ �p��[-�k���f���R�D!��Z#��D!��T
%)�u:=�o7���x�n�����l����]�w;����Z������L�c1,���~�@  0���O'��B��@��P$29.�[-��u�}>?���s��N����H�b��R�D�a�x.7�M&3�L�c����C!����E�q�|����z��G#�r��F��`(�z�N�C�P�d)��U�u:�^���p,6�].�[�V�E"������p,�{������|�o7#��R	�b��Y,6;�����x.7�M��y<>��o7��C!�h��z�g3�s9.��m�{=�o��m�{=��k5��v�M��y<>?�C!�h��U*�Z�F  08<��_�W+�e2���G#$2�\'��d�T
���d)�j���b$�y<��_�W�U�u:��O'��d��J!�h*�Z�F �p�v�M&��l+�����h*5�����v�M&�Y�v�M�s9��{=���{���g3��F�A��X��S����b$2�\'�����d)*5��v�M�s���G�Q(���n�P�r�f�I���������l+�e�y��_�W+
�R	�b��D�a�x�n�B  08�~�O'	�b�d�T�e29���k���f�I���l�U�u��~�@�`(����W+
%)�j�J!(�z'�I$���^�G#�r&3�s9.7�M&����K����R�D�a0�|�o��m6��n�E"1,6;�S)�u��~��g3�f��B�`�t��v#�d�i�z'�I���l�k5������[�V�B�`����E"�X&3�f���A 0��^  �x����u�}>?����X�f���R��B����D�P���l��j���b��R	"1�l+�J!��T��r�L#�H"�X&3�L#��R��B�@�`��T�e29�n����Y��[-����]��{�^�`��T��r�s9��W+��E�q8<>�_/���r��F�`�h*�Z�F��������`�h*5��v��C�P�d)�u:=/�B ��X��y��_/�a��\'�I$29���k5�V��b�r�L��q�|��w;���c��L����J�P���I�r��F�A�p���K%���Z#��Y,��}>?���s9�n��������b���B��@�`(�z�g�Y�v�M�����O'	"�X&3���C!�h�u��~���s9.�[-+�e2�\���t�V�������E"1,��}>�_/��e29�n�����l�k�Z���T��r������M�s���G#$��|�����~��P��R	�q8��_��k5-�k����S)*���f�I�r����^�C!�t��K%)���j�J�����A 0�|�W���U�u:=�W+��r&��l�k�Z�F��`�t�V��A 08<>?���p�v��q8<>����{��O'��d�i4�}���o�[-+
���d���Z�F�A 08<�?��c�X��S)�u��~��g3�L#��D�a08�����{=�o����[-��j
��I$����O�S)�j�e29.7�c��L#$�y�~��g3��������F���@�`(4:=��w;������O�S)*�Z�F��`�t���[-��u:��O�S)�j���Y�v�M&��l+���Y�v�M&3������M������g��l�k�Z�F��@ ���L��q�|/���r�L�Q�t-�k����S�T������K�R�D��p�v�M&3����a0�|����}>?�O�S���E�q8��_/��A �x�����z�S�T��r&��l��j�J���X&3���C!(4:=/��A �����c1,6;�N��`�h�j����Q(�����k��M���|����}����?�C�P$29�w;���t-��u:=/�K%��t-�k����S�T
�R	�q��^�G#�d�����Q(�z'��B �p��V����h�u:=�o��m6���W+���b�d�T
%�i4�}��?�G�����E"1���K�����I$�y<>�_/�B�@ �p��V�E"1�l��j
��I$29.���v�c�X&3&3&�Y,�{=�o�[-�U*������t��v�F��`(�z�N��a08�~�O'�I$29�n�E�q8�~�G��h*5���[-+��r����t���[��K�R	�b�H��Q(����W+
%�T�e���^����H"�X&3��F���P$2�\'	�q�|�o7��q�|��w;���y<����_�W��j���Y����v������G#�H"1,��}�?��g�����e2�\'	"1��V��b�d���E"1��V!(4:=�o7�F�A��X��S�T
%�i��].7��h�j
%��t��K%�����f��B��@ ��X��S�T
%�i4:=���u��~��c���F�A��X�s�\�S���E��x�n��e29.7������Z#��D����L�Q(4:�^�G#�H"1,6;�N��a0�|����z����|�o��m6�]��{�^����x.7�M&3��F�@��P$�y���o7�����X&��l+��r&3�f���R	"�X�f�D!��Z#�H��Q���M&�Y��[-����j�e��|/���Q�t�m6;�g3�s9�n��b$�y<���_���u�}�?��g���V�B��P���l+��E�����G�Q�t����m�{=/����Y�v�F�`�t�V���Q�t-+��E"1��V��p,6�]�w�]�w�].7��q8�~�O�S�T�e��|��k�Z��q���O���t�m�������{=�W�U*5��v��q8<�?���q�|��k��M���|��w;��G#��������D!�h�j
%�T
�����I�r�L�c1�v�c1�v�M&�Y,�{=�W�U����n�K%�T
���d�i������u�}>?�������A��X&3�L#�d��J�B��������P$��|�o7��f�D�����F�@�`��T
%�i4�}>?�C��H��x���k5�����Y,�{�^��c�X����^��c��L���x���k�Z�c�X�f�����P�r���i�z��i4:=��w�]����~�O�S)��U*�Z��q8<������}���_��k�Z#$�y<����_�W�U����n�E�q8��_�W�U*�Z�F��`(4�}�����w;��i�z�N���p�v����\��s����c�X�f	�b����V�B  �x��{���g��l�k5�V�B  ��\�g��l��u:=��w;���c1�l�k5����r�f�I$�y�~��c1�v�F���@����D�P�r��S)*5-+�e2���G#�H�b��D!(4:�^���q�|/�K�R	"1��V���������Q��Z�F  0�|�o�[�����Y,�{�^��`�h��U�u��~�@  0�|/�P$29���}>�_/�K��I�r&3��F���P�r�L#�d��J���D�a��\'�I���l�k�Z#�d�i����W+
%��t�m6;�S�T�e29�n�K%�i4:=�o�[��K%)�u�}�?�C��H"1��[-+��E�q��^�C!�h���]�w�]���}>�_/��e29��W�U��z��s9.�[-��u�}>����{��O'	�b��R�D���D����B�@ ��X&����K%)�j�J�������a��\'��B  08<>�_�W+
%�T
��I$��|��k��M���|�o����[�V���Q(��]�w�]�w;�N�����L��q8<>����{��O�S)����n��b�r��F�A ��\'	"1������Y�v�M&���V�a��\��i4:�^�G�Q��Z#�H��������x��{=/���r�L�c1,�{=/��e�y<>?�O��i��].7�M&�Y,6�]�w;�N��`���������M&��l�����n����Y,6��n��b�d)*5�m6�����u�}>������~��g���V������J�����H"1,6��n��e29�n�K%)�j
�R�D���X�s���G�Q�t�m��}>���w��n�K%�T
���d�i�z����������q8�~�O������f�I$2��N��`�h�j
%��J�a�x�n��e�y����w;��s�\'�D!�h�u:���g����K%)���].�[�V�E�q8<��?�G#����A 0�|/��b���I�r��F�A �x���k���f����I$29.7������L#��Y,�{����s�\�g�Y���m6�]��{�^�A ��\���y�~��c���F��P�d)����n��e2�\��i4:�^��@ �p������Y,��}>?��a0�|�o7���a����G#$��|�W+
���d�i4:��O�S������h�j���b���I$2��N��@ ��X���i�z�g3�����p�v���x.7�����t�m6�������].�[���e29����u:=/�E"1,6���W+�J�a08<���_�W+�J�a�x�n��p,����_�W�U����n��e29���}�?���p������Y,������w;�N���p,��}�?���s�\��s9�w;����|�W+���Y,�{�����y<>?��a��\�S��J!(4:=�W�U�u�}>?�G�Q(4:=/��b�H���h����U�u:�^�`(4�}>��o���v�M&�Y��[�V���D�a0��^�A�p�l�k5�V��b�d�T
%)*5������[-+
%��t�V���Q(4���_/��b�����`�t���[�V�E"�X&�Y,6;�������S����b�d��t�m�{�^��a��\'�D��p�l�k5�������m��}>?�������O'�I$��|�o�[-����j�J�B�@  0��^��a0��^�G#�H��Q��Z�c1,6��n�K%)�j��r�f�I$����O'�I��Y,�{=��w;����|��w�]�w;�N  08<>�_/�E�q��^�C�P$���^�@  0�|��w;�N�A�p�������l+��E"�X&�Y���m�{=/�K%�i�z����q�|���{=/�E"��L��q�|���u�}�?���q�|�o�[�V��A 08�~�O'�I$29�����z'�D!���J��A�p������Y,���~��g��l+����Q(�z��s�\'��d)*��M�s��N��a��\�g3&3�L��q���O'�D�P�����K%�i4��~�G�����E"�������X�����Z�c�X�s9��W+�J�a�x�n���Q�t-�����n��b$���^��a0�|��w��n��e2�\��s9.7�M&�Y��[-���z�����^�G#�r�f��d��t-��u:��O'�I�r���C!��T
%���E�q��^�G��h����U�u:�^�G�Q���M��y����w;����q�|����}>�_/�E�q�|��w����k5-�k5-+���b�����`�h��z����Z�F�A ��\�g3����a0�|�o�����m�{�^��c1�l�k���f	��Q(�z���c���F���@ ��X�f�����P���l�k��M&���V�E"1��[-��j�J��H"1��V���Q�����S����b���B��P�d��t-�U����n��e��|���u:�^�A 08�~��a�x���k5�m6;�g�Y�v��������f���A�p�l�k���f��d�i4:=/�E��x�����z���y<��_/�B�@  08<��_/����Y���m6;����Z�F�A�p�v�F�@�`���M��y<>?�A ��\'��B �p,��}>?��g�Y,��}>�_/�����T
%����M��y�~���P��Y,�{=/�K�R��������B�`(4:�����y<���?�O'�I��Y,�{��O'�D��H"1���K%���Z��q�|/�K����R	�b�d)�j
��I��Y���m6�].7�M&3���i4:=/��b��R	"�X&��l��u��~�G�Q��Z����p�l�U*5��K%�T
%����M&���V��A�p,�{=�o��m�{=�W+��r������X&�Y�v�F�A �x��{=���{=���u�}�������w���W��j�e2��N���p,6���W��j�e��|/�E"1��[����r�s9.7�M�s�\�g�Y��[�V����P$2�\��i�z���y<>?��`����f	���\���t��v#�d)�j
%���Z#��R	"1�v�M�s���G#�H���h����n�K%�i4�}>��o��m6������z����q8<>?��g���V�P�r��F�A �x��W�U*5�m���~��g3�L�c1�v�M��y������}��?��c�X�f���A���L��q8�~�G����J��A�����C������`��T��r��F�A��X&3��y��_/���r�L�Q�t�m�{=��w�].7#�r�L�c����C!����E�q�|��w�]���}������w;�g3����a08�~�G#�d���E��x�����z�g�Y,6;�g3���C�P�r�f�I����V�E"1��V�E"1���m6�]��{=��k5����m6���W�U��z�N �p��V�B�������`�h�u�}>?��g���V���`��T
�R	��x���}>?�G��������h*���f��B  ������q�|��k5��v���a08�~��g3��F��@�`(4:=���{=�o7��f�D�a0�|�W��j
�R	��x�n�E�����G#��D����L#�d)�j�J�B�@ �p���K����R	��Q�t��v����i����W��j�J��A��X��S)�u:=�W�U�u:=���u:=�o7��f	"��L���x�n����h�j
��I�r�L�c�X�f�I���l�U*5-+�e2�\�g�Y,��}�?�����\'���R	�b���B�@  08��_/���Q(4:=��w;�g3���C����B  �x�n�a�x�n������C��H�����J�P$29�n���r�L�Q�t��K%�T�e29��{�^�G������b$�y�~����x�w;����|�W+�J�a�x�n�K�R	�����J��p,�{����s9���k5-�k5�V������D��H�b��R	�b�H�b�H"��L������G���T
��I$29�w���W�U*5��v�M�s����c�X�f	"1��V�E"��L������b�d��J�B �p�v�F �����C!����f���A ��\���y<>?�O'��d���E��x��W+�e����O'���R	���h�j�J�a�x.7#��D���X��S)���j�����V��b�d�i4:�^�A��X&��l���z��G�Q�t�m6����k������t���[-+
��I$��|����z���c1�v�M�s���G�Q(4���_/�K%)*��M&������r&�Y��[-�U*5����r�f�I$29���k�Z#���B��P���l+��r���i�z��s9��W�U*��M&3��y�~�O����Z�F�A�����C��H"�X��S�T
�R��B ���L#��Y,���~�G#�d��t�V�E�����G#��D��p,6�].�[�V���Q(4��~�O'	�b�d���Z�F�A 0��^��a08<>?�A 0������y����w�].7���S�T
�R	�q8�~���q��^����X���i4:���g��l��j��E��x�n�K%�T
�R	����T
%���Z����J������D!(����W+�J���D���X�f���R	"1,�{��O'���R	�q��^�G�Q(4:=�o�[���e29�n�E���������\'�D!��T��r�f�D�P���l��j
�R������H�����G#�d)*�Z��q�|�o����[�V�E"1�v�M&3��y�~�`�t�m���~�O'���R	"1�l�k�Z�c1��V�B��@ �p�v#$��|/�K�R	"1,6�]�����_�W�U�u:=/���r�s����c1��V���Q�t���e�y<>?�O�S)�j
%�i���n��A 08�~�O�����M�s9�n�K���d�i4:=�o7��h���]��{=���{���g��l��u��~�O�S)�j�����V����P�d���Z�c�X�����Z�Q(��].7��f����I���l�k����S)��U*�Z����p,�{=�o���v���S�T
��I$29�w��n����P�d�T���Y�v�F�A 0�|/�K�R	�q��^�G��h�j����Q(4�}>����{��O�S)��z�N�C�P����V�a0�|�W�U*��M&��l��u�}�����o�[��K��I$2�\��s���G�Q(4�}>?�O'	"���F �p����e��|��w�]���}>���w�].7�M&3���C!����f�I$�y<>������~�O�S��J��A �x.��m�{�^���p�v�F�A 0��^����D�P����d������S�T
%��J��A �x��W���U*5-�k�Z�F�@�`�h*5�m�{=���{���g3��F�@ �p���K%�i4:=�W��j��r�s9�w;�S��J���`�h�j�J�a0�|�o�[-+
%)���j
�R	��x.�[���e29��{�^ �p�l+�J����P$��|�o7��f�I��Y,���~�O'����I�r���|�o7#���l�k5-+�����V�P$2�\���y<����_��k��M&���V�����T
%)�j�e�y<>�_���u:��O�����M�s�\��s9.7����i4:�^���p,6�]�w��n�E"1�l���U�u:=�o7��h��U�u:=�W+��E"1���K%�i4:��O��i�z�N�C�P$29.����[-�k5-�k�Z�c��L��q8<�?�O'�D���X��y<>�_��k5-�U�u:=�o7��f���R�D���X�f�����d��t-�k5��v�M&3�L�c�X���i�z�����x�n����P�d�i���n�E"1,6;�S                                                ��G                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   �         ��          �                                                                                                                                                                 �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    ��    ��    ��    � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���������������������������������   � �� �   � �� �   � �� �   � �� p   � �� x   � �� `   � �� h   � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��      � ��         ��         �� �      �  �      �                                                                              ����  ��������������������������� ����������������� ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                �                                                                                                                                                                                                                                                                                                                                                             @                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        