1VSB    $�8ё> BST1   $�8�Compatibility                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �   ��@� ��@� ���b    � 7 ��  6�    �� ��ߤ�                      ]    ��  @�����@K K               � �                                                                                              p ��  
   �'R)�)R+�)R+�R�!R#�zR|                      � � ��                                                                                     �         @                                                                 ^ � 6o  ^ � o  f � o  f �  o  V � o  V � o  U � o p m   h m  " p &m   � +m    � +m  " h  m v .m �� b* �� d* �� d*   ��  + �� +   �� +   �� +   �� +   �� +   �� +   ��  c   �� )  � {  j � � j � � j � � j  � � j  � � 
j  �� c   �� c  � � b*� � b*  � � d*��n i  ��f i   n &i  ��� +i    � +i   f  i��t .i d c   \ c   d &c   z +c   z +c   \  c j .c$ a a  $ Y a  , a &a  % w +a  * w +a  , Y  a# g .aH a e  H Y e  P a &e  I w +e  N w +e  P Y  eG g .ed g g  d _ g  l g &g  e } +g  j } +g  l _  gc m .g �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �       �      ���9��  ���=��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ^�6o^�of�of� oV�oV�oU�oomgm"o&m�+m �+m"g mu.m�z j��j��j��j��j��
j�b*�b*��d*�mi�eim&i��+i �+ie i�s.icc[cc&cy+cy+c[ ci.c$`a$Xa,`&a%v+a*v+a,X a#f.aH`eHXeP`&eIv+eNv+ePX eGf.edfgd^glf&ge|+gj|+gl^ gcl.g��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��         ��b�� ( 
                                                                                                                       p    � X  ���������������������������������������������������������������������������������������������������������������� ��� ���!���"���"���#���#���#���$���$���%���%���&���'���'���(�������������������������������������������������������������������������������V�V��������uMlM|MuM#M - -(181H1X1e1;1�����������V�V���������ul|# - -)191I1Y1K1[1=��=��>��>��?��?��?��@��@��A��A��B��B��C��C��C��e *�d *�d *�d -�d 0�c 3�c 3�c 6�c 9�c 9�b <�b <�a ?�a ?�a B�a E�a E�` H�` K�����                                                                
                                                                                        ��W ��W ��W ��V ��V ��V ��V ��V ��U ��U ��U ��U ��U ��U ��T ��T  �O`��T ��T ��T ��S ��S ��S ��S ��S ��S ��R ��R ��R ��R ��R ��R `   `   `   `   `   `   `   `   ��P ��P ��P ��O ��O ��O ��O ��O ��O ��N �� I�X  �  ��  �  &1 *  �X �   ��  �B �@ 0+DQ"S*"R2#���� �� �$ � �. 8* 8. 8, 8( 8" 8  8$ 8& &1� � � �� =� M� 6� Q  /K (Z C8 2 7T =Y     �,�  � B� �G & 2# F � � � ,� *� � �� ��   �  �  d  D  V  n  �  �� �4 �O �� �� �� � �) �& � # � � � Z� \  ?�J' \ � � �X��I! IJ�;0R ��@�@��C��C��E ��  � �� @� �| @{ @{ ���[�6��7��9��;��>
���պ �� ׷ �� �� �� �P ��     �P                                                                 ��  ��  ��  �   �   �       �� �m an 9� j* j* �� �n {" �F 2;                       	  	  	                       ��  ��  ��                                         a                                          -�- -8-(-`-�-�-     	  	                                                                                                 �  �  �  �  �  �  �  �   �   �   �   �   �   �   �   � �    �   �   �   �   �   �   �   �   �   �   �   �   �   � �Y� � � �  �  �  �  �  �  �  �u��5�U��x�`�$�T�.��t�%�z�v�}����/�!�?�6��9��J�<�|�W�-�y  @ �b�c�d�=�,�f�e�g��4�I�r�hiO|q{jx[xVvpukt>s3rHpooln]mkjn  @   @   @   @   @   @   @   @ UEMsMM&IKG*F^FE+DDB<<M<';_;:1:F:6C4L/,D,@)~){!G A                                             ������
                                                                                        � �                                                             � � U �  i ��g  ] # Z G Z c `                                                                   ��                                                              ��  ��  ��  ��  ��  ��  ��  ��                                                                                                                                                                                                                                                                                  � �  �  �  �  �  �  �                                                                                                                                                              �k��          C[  �                                                                       
   
                                                                     �  �  �  �  �  �  �  �  �                                                             ��  s�  ��  {�  ��  ��  ��  ��                                                                  U  �     �   �  �  �                                                                                                                                                                                                                                                              ��                                                             @  �������_���q���������������                                                                                                ��                                                            ����l�L�^�v�����                                                                                                                                                                                                                         �����  �  0 X                                                                                                                                                                                                                                                                                                                                                                                                                                                                 l                            �_�g�1�-�6�W��%2[�  �%O�HA�!v!�!�-�6�W�1W6=S�w�!���#9g��yu�{����(�)�)d*�#�H1'e0S�[�g�g�R�c�k�s�{����#9g�Y9YB�J9K;�Q�Z�s�Q)�5_[�#��9�#�#�#�G��{���S�c�s��-9g�S9WB�J7K�1;�Q�������#9g�T]Xfg8g�1_�Q��0S�_�o�{�:     �� Fp ?'W�k�_Q  �AU=�$�eF �U�~?W�k��G  � e ��F �?W�k�k  �E� hb�F q�_?W�k�9~  
E$ qe�8F �}_a?W�k��  � �� F�?_'W�k��  nD%��iNF_!Ng?'W�k��1  B$�$ �@�8F k]_Q?W�k����� �UU @33�*�$  q�EU�I 8y�0�!�
=
�	{	$	��B ��P���f>����rU9�����}iVD2! ���������ui^SH=3)�����������������|vpjd^YSNIC>940+&" ������������������������������������������}zxvtrpnljhfdb`^\ZXWUSQPNLJIGFDBA?><;9865320/.,+)('%$#! 
	 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ^�B                                                                                                                                                                                                                                                                                                                                                                          ��                                                                                            ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          �)                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ��������������������������������������������������������������������������������������������������������������������������������:     �� Fp ?'W�k�_Q  �AU=�$�eF �U�~?W�k��G  � e ��F �?W�k�k  �E� hb�F q�_?W�k�9~  
E$ qe�8F �}_a?W�k��  � �� F�?_'W�k��  nD%��iNF_!Ng?'W�k��1  B$�$ �@�8F k]_Q?W�k�  �_�g�1�-�6�W��%2[�  �%O�HA�!v!�!�-�6�W�1W6=S�w�!���#9g��yu�{����(�)�)d*�#�H1'e0S�[�g�g�R�c�k�s�{����#9g�Y9YB�J9K;�Q�Z�s�Q)�5_[�#��9�#�#�#�G��{���S�c�s��-9g�S9WB�J7K�1;�Q�������#9g�T]Xfg8g�1_�Q��0S�_�o�{�:     �� Fp ?'W�k�_Q  �AU=�$�eF �U�~?W�k��G  � e ��F �?W�k�k  �E� hb�F q�_?W�k�9~  
E$ qe�8F �}_a?W�k��  � �� F�?_'W�k��  nD%��iNF_!Ng?'W�k��1  B$�$ �@�8F k]_Q?W�k�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  l-l/                                                                                                                                                                                                                                                                                                                                                                                                                                    ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                                                                                                                                                                                                                                                                                                                    �������������������������������������������������������KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;� � � � � � � � � � � � � � � 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�{�0�{�0�{�0�{�0�{�0�{�0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      # ���       �      + P               �Q                                                                                                                                    �� ���������
������                              �����������������                              ��� ��
���!���
�
�!�"���                              
�
�#�$�
�
�
�
�
��
�
�
�
��
�
�                              
�
�
�
�
�
�
�
�
�
�
�%�
�
�
�
�
�                              
�
�
�
�&�'�(�
�
�)�*�+�
�,�
�
�
�                              
�&�'�(�-�.�/�
�0�1�2�3�
�4�5�6�
�                              7�-�.�/�8�9�:�;�<�=�>�?�@�A�B�C�7�                              D�8�9�:�E�F�G�H�I�J�G�K�L�M�N�O�D�                              P�Q�R�S�T�U�V�W�S�T�U�V�W�X�S�Y�P�                              8�9�:�;�<�8�8�8�8�8�=�>�?�8�@�8�8�                              A�B�C�D�E�8�F�G�H�I�J�K�L�M�N�8�A�                              O�P�Q�R�S�T�U�E�V�W�X�Y�Z�[�\�]�O�                              ^�Q�Q�Q�R�S�E�_�Q�`�a�b�Q�Q�c�d�^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                � � � �B�a�a�Q�Q� � � � � � �<�b� � � � � � �!�A� � � ������ � � � � � ���� � � � � � ���&� � � � ��@���(� � � � � � ���L� � � � � �p����� � � � � � �� � � � � � � ���@� � � � � � ���L� � � � � � �8�E� � � � � � ���� � � � � � � � � � � � � � � � �I�I�E�C� � � � �A�A�#�� � � � �I�I�[�6� � � � ����� � � � ���6��� � � � ����!������ �h������ �`��� �D�D�D�B� � � � �x����x� � � � ���	�� � � � �@�����`� � � � �D�D�D�B� � � � �������x� � � � �$�$�l��� � � � � � � � � � � � � � � � � � � � � � � � � � ��� � � ����9�f� � � � � ��B�b� � � � � � ��"� � � � � � ���L� � � � �� ��� � � � � � � ����� � � � � � ���d� � � � � � �p��� � � ����?�� � � � � � �<�b� � � � � � �\�2� � � � ����� � � ������� � � � � � ���$� � � � � � ���@�:�D�N�;� � � � �B�B�F�;� � � � �$�4��� � � � �~�@�b�<� � � � �D�D�D�B� � � � � � �2�� � � � �������z� � � � �E�A�A�@� � � � ��� ����� � � � ����� � � � �A�A�#�� � � � �"� � � � � � � ����� � � � ���$��� � � � �/�H�L�'� � � � ��� �@��� � � � � � � �A�C�&��� � � � � � �<�b� � � � � �8�D�`� � � �@� � �.�1� � � � � � �A�B� � � � � ����,� � � � � � ��� � � � � � � �8�� � � � � � ���L� � � ����r��� � � ������ � � � � � ��� � � � ������F� � � � � � ���$� � � � � � � � � � � � � � � � ����� � � � �A�A�#�� � � � �<��B�<� � � � �!�"�"�!� � � � �G�D�f�3� � � � ��� �(��� � � � �����@��� � � � �t�����v� � � � �D�D�D�B� � � � �������v� � � � ����� � � � �'�(�i��� � � � �D�����k� � � � �$�"�b������ �@�@����� � � � � � � � � � � � � � � � �!�s�U�I� � � � � � ��� � � � � � �\�2� � � � �@� ����� � � � � � ���@� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �A�A�A�!� � � � �:�D�N�;� � � � �"� � � � � � � �������c� � � � � � �`���� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�+++��++++�+++�+����++�++++�+++�+��++�������+�+���������+�������������������+�������������������������������������������D�D������DD�D�D����D�D��D�����D�D�����DD�D�A�AD�D���D�D��D�D�A�AD�D���D�D�����A�A�A�A���A�A������A���A�A�A�A���A�A������A����A��A���A�����+������A��A���A�����+���A�++++�+++�+�++�A��++++�+++�+�++�A�����������������������������������������������������������������������������������������������������������������������������������������������������������������*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�j�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�j�j�*�*�*�*�*�*�*�j�*�*�*�*�*�*�*�*�j�*�*�*�*�*�*�*�*�*�*�*�j�j�j�j�ꢪ*�*�*�j�j�*�*�*�*�*�*�j�j�j�*�*�*�*�*�*�*�*�*�*�j�j�*����*��*���*�*�j�j�*�*�*�*�*�j�j�j�j�*�*�*�*�*�*�*�*�*�j�j�j�*�*�j�*�*�*�*�j�*�����*�*�*�j�j�j�j�j�*�*�*�*�*�*�*�*�*�j���*�*�j쪢����*�j�*�j��j�*�*�����j�j�8�8�8�*�*���*�*�*�j�*������*�*�j�*�*�*�j�j�*�*�j���*�*�*�j��j�8�8쪈���*�j�*�j�j�*�j�j���8�*�j��誢j�*���*�*�j��j�*�*�*������8�*�*���j�*�*�j�j�*��j�j�8�8�8�*�*�j�*�*�ꈪ�*����8�*�*�*�j�j�8�*�*�*�j�j�*��j�8�*�j�8�8�8�8�*�j�j�*�*�j�*�*�j���8�8�*�*�j�8�8�8�*�*�j�8�*�*���8�8�8�8�8�8�8�8�8�8�8�8�*�*�*�j�j�8�8�8�8�8�8�8�8�8�8�8�8�*�*�j�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8sss s�8???�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8{{{�x�x�x�x&s$s"s@s ?"?$?&?�8�8�8�8�8�8�x�x�x�x�x+++�8�8�8&{${"{ {�x333�8Bs`s@?B?�8�8�8�8�8�8�8�8sss�x 3"+$+&+�8�8�8�8�xB{@{ 3"3$3&3�8�8s`3333�8�8�8�8�8�8&s$s"s s@3B3�x�x�8kkk�8�x`s@3B3�8�8�8�8s(3"3$3&3�������X�xBs@s`3�x�X�X�&k$k
;;;s`3��{{{({H3B3�����������X`sJ?L?� ;";,;&;D3F33�8&{${"{H{h3������������x{j?l?&$" @?B?`s(3d3f3&3�8�8�8B{hsJ?L?�����ssssj3???B@`3�sH3b3N3{{�8�8�8FsDsl?&$" �;;;&s$s"s(s(?"?$?&?�`sJ?L?s`3sn3${
???{fsds s��B@ ;";$;&;��BsHsH?B?��LsJsj?l?s3sJ?L?"?$?&?&{ 81          � � � �����  � � ` ``� �    <=              � � � H����    � � p  00�0          x              8         � x�4��          ` 8    8|6�>�>��   6>>wl` � < :$rL��✁�   @ �$�L�� �@�  !@?@?�I�I�I�            � � ����ܸ�|�  � | p ��������  / � �          /   @ � � � � � � �     � � � � �  � � � � � � � � � � � � � � � �     � � � � � �       �    2                                   $(	
	
         ! 8<          \����0�� � � 0�`�� � �   sC<A>8   3       ������0�� �� � 0�� � �   |���~�b@ > < y s  ?    ������|�� � �� �� �   I9�g�ow?  9go       ��b���� |�� � � b�� �   �     �~?|7!> 8? ??77      |�� � � < ~  � ��x X � � � �   |� o �/  0 0          ���� 80��� @ �8 � � �                          p�p �          P                ~ �~�~�             ~  � � � | ?      ` p 8       /+/'          � 0�� � Ԁt ��   @ � � x � � �   @&@ �H�@                � 0�0                      @&�F�P                    � �                                    �  �                   9yk�0�0�     0 " F O  � � ������  � � � � � � �                                        � � �             � �  @#@'@'�O�O�O�G               � � � � � �                     $f$�Z�[f$$ < ~ ��$�$�~ <      <<          < <      ?:/.              ��(�H���0��� � � � � � �     �@�@@ @                   "$00��                �@�@@                       "$��                                        $(HP  ��        @        � �  @     o O 0 ?       ��<8����� p 0 � � �       >>               � � � � � 0 �08 � @ x � ` �            $                     < ^ f f z<                      <f$f$<      < ff<                                 �������G  < | ~ ~ ~ | 8 � �������    < < <  3gN1�"�@�@      � 8��0�����       ����������� � � � � � � �          � � � � � � � �   � � � � � � �     ` �`�p�pL0J4                 $$&I6I6�l�                         ?                   � � � � � �                  <B=�x�p�c`'p        @ � ��0���     � �p0p  @8`0p�;�           � ��,��      � �00�p �p�xa@?I68                 ` �`�`H0H0�x�\a                ���x�p�p�p�?       O@08   ���~~y~�� <   ���x�   �@�p�0O0o0           � �3��<0��� ������ 0��   !!    ��!!    ��� � � � � � � �     @ ` � � � � R,B<F8I6�~�l�``                 		`�|�nn                 ?    � � � �                 � � � � � � � �                 �~�|�~�L48  @@` 4   ���np�� p ��  ��| � p  �~�~�N>6  @` >    |��s|Gx>�� � �� ��~�~ � �        � ���p�                  ���p�x�l�ny                                                                              ~~����~~xx��cc  ~ � � ~ x � c77������   7  � � � ���������������� � � � � � � � �00yy{{kk    0 y { k �����������ޞ� � � �  � � � �      00            0             ��          �   qr���p�``    0 d h        0@0�c�g�           @� x�$���      � �8� 9 %"0            � �\���pp ����    � � p� @ @ ? oP?W8T8W8_?`         � ����8T8�8���  � �    � �   <<~~~~<<  ��     < ~ ~ <   �    <<  @@      <    @     ll������8888   l � � � 8 8 ������?????? � � �  ? ? ? ���������������� � � � � � � � �����qq##99 � � q #  9  TT����^^LL����   T � � ^ L � �      !!           !        ��  ��      �     �    < B<�v�b�B�fB<<                 �~` `?r>_?# `    2 ?   ~~��4848�� ��� ��8�8 �               ��������� H  � @ @ @ @   ����  ?            � @�x�h�x�h�H��   � � � � � �                                                                                                                                                      �? � � � � g             � � �� � � � � �              @ � �o�m�#�#@    0         �����@�������p� | 0        � ��������v���              �ց��ԃԃ����� � ( x ( ( 0     ? � ����@?@?@?           � �� ������ � �           #�?@�`� � ��g�             |�� � � ���`             @ �  ` �`��d�| �           �                                                                                                                                                                   � h             o               	 �   � � �       L0�|� � � � � �          0 �     �p� � ~ <�{�1� p     � �    � B�<��( ��<~ <    � �   �p� � � ���� p         � � � � � � � �                 � � � � � � � �                C Q ) &�"���� � � � A A a    � � � { 3   �        � � � � 7 � � � � � �               p � � �          ��          ��          ��          ��          ��          ��                              �          ��          ��          ��          ��          ��          ��                              �          ��          ��          ��          ��          ��          ��                              �          ��          ��          ��          ��          ��          ��                              �          ��          ��          ��          ��          ��          ��                              �          ��          ��          ��          ��          ��          ��                             �s�s�s�s�s�s  ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������       �Z�N��G        ��~    @   �B         Da~   ~ � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � dfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLN      
    
             " $ & ( * , . 0 2 4 6 8 : < > @ B D F H J L N P R T V X Z \ ^ ` b d f h j l n p r t v x z | ~ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �  
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPR      
             " $ & ( * , . 0 2 4 6 8 : < > @ B D F H J L N P R T V X Z \ ^ ` b d f h j l n p r t v x z | ~ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �  
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`bdfhjlnprtvxz|~���������������������������������������������������������������� 
 "$&(*,.02468:<>@BDFHJLNPR      
             " $ & ( * , . 0 2 4 6 8 : < > @ B D F H J L N P R T V X Z \ ^ ` b d f h j l n p r t v x z | ~ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �  
 "$&(*,.02468:<>@BDFHJLNPRTVXZ\^`b�  ~ H * � ��@  #   �   ����X�X�X�      �    K   K                                                        l  l                       @                                                                                                      U���@���\ �~\��~@UUUUUUU9  K           =                                            UUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU ��� B   ���   �   0  �ް�    %".�   �         �   P   �                                                                                                                                                                                                                                       ��        ��        ��        ��        ��        ��                                                                                             ,                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        ��������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������                                                                                                                                 � � � � � � � � �                    � � � � � � � � �                                                                                                             ��0                 ih:4w     "     ,U~^8p�@P~5p  @P~5p                                                                                                        ��                                                                                                                                                                                                                                                                                                                                                                                            �                        �X�Z�\�^                                                                                                                                                                                                                                                                                                                                                                                                   `6                                                                                                                          ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              z     @ 	
@ABCDEFGHIJKLMNO 	
@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_PQRSTUVWXYZ[\]^_ !"#$%&'()*+,-./`abcdefghijklmno !"#$%&'()*+,-./`abcdefghijklmno0123456789:;<=>?pqrstuvwxyz{|}~0123456789:;<=>?pqrstuvwxyz{|}~                                       �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	
		









		
	
	
 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~��������������������������������������������������������������� 	
 !"#$%&'()*+,-./01     ! " # $ % & ' (***************888888888888 >>>>>>>>>	>
>>>>>>>>>>>>>>>>>>>>>> >!>">#>$>%>&>'>(>)>*>+>,>->.>/>0>1>2>3>4>5>6>7>8>9>:>;><>=>>>?>;;;;;;;;;;;;;;;????	?@ABCDEFGHIJKLMNOPQRSSTUUVWWXYYZ[[[[\]]] ^ iiiiiiiii	i
iiiiiiiiiijjjjjjjjjjjjjjkkkkl�	�
������ �� �� �� ������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  � �����-�-�-�-�-�-�-�m�6 �- *****
***�m�6 �- *"*$*&*(***,*.*�m�6 �-@*B*D*F*H*J*L*N*�m�6 �-`*b*d*f*h*j*l*n*�m7 ���������������������� @ABCDEFGHIJKLMNO��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        H`6��{~�H�}� *p� H�~� ,p� &H�� .p� 2H�� .p� >H�
  ��_  JH   ��_  VH�  ��_  bH    �_  nH�   �_  zH   @�_  �H�  `�_  �H   ��_  �H�  ��_  �H   ��_  �H�  ��_  �H    �_  �H�   �_  �H   @�_  �H�  `�_  �H   ��_  �H�  ��_  
I   ��_  I�  ��_  "I    �_  .I�   �_  :I   @�_  FI�  `�_  RI   ��_  ^I�  ��_  jI   ��_  vI�  ��_  �I 0�
  �I  � (p �I                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������A��A��B��B��C��C��C��e *�d *�d *�d -�d 0�c 3�c 3�c 6�c 9�c 9�b <�b <�a ?�a ?�a B�a E�a E�` H�` K�` K�` K�_ N�_ N�_ Q�_ T�_ T�^ W�^ Z�^ Z�^ Z�^ Z�] ]�] `�] `�] c�\ f�\ f�\ i�\ i�\ i�[ l�[ l�[ o�[ o�[ r�Z u�Z u�Z x�Z x�Y {�Y {�Y {�Y ~�Y ~�X ��X ��X ��X ��X ��W ��W ��W ��W ��W ��W ��V ��V ��V ��V ��V ��U ��U ��U ��U ��U ��U ��T ��T ��T ��T ��T ��T ��S ��S ��S ��S ��S ��S ��R ��R ��R ��R ��R ��R ��Q ��Q ��Q ��Q ��P ��P ��P ��P ��P ��P ��P ��O ��O ��O ��O ��O ��O ��N ��&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&�&&�&&�&&�&&&&_&&?&&&&�&&�&&�&&�&&&&_&&?&&&&&&?&&_&&&&�&&�&&�&&�&&&&?&&_&&&&�&&�&&�&&�&&�&&�&&�&&�&&�&&�&&�&&�&&�&&�&&��������������������������������������������������������KKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKKK;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;;� � � � � � � � � � � � � � � 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�{�0�{�0�{�0�{�0�{�0�{�0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� 0�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � vAj  ,�Z~pp C]~_A �	�	�                                                                                                 pp C]~_A �	�	�	�	�	�	                                                                                                 ��V�tX C�[~� R� R C!\~ "\��S                                                                                                 �,U��U C!\~ "\��S"\ &&�C\~                                                                                                 �@P�Q C�\~ �U��U�U A&�\~�U�                                                                                                 �U��U��V  Z~vj  ,�Z~pp C                                                                                                 _A �	�	�	�	�	�	�	�	9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ���++++�+++�+����++�++++�+++�+��++�������+�+���������+�������������������+�������������������������������������������D�D������DD�D�D����D�D��D�����D�D�����DD�D�A�AD�D���D�D��D�D�A�AD�D���D�D�����A�A�A�A���A�A������A���A�A�A�A���A�A������A              ?         ��������        ����3��        ��89899        ��?���?        ��������       �?8��������        ?       |��������   ""D������ݻ;   ?  `|�����ߟ�   ��������   8��������  <FBD$��ù����     !A������޾���37?ll�����    ��������s!,                 �         �        ��������        ��      ��������0@�   �Ͽ�����x  ����3���Ƅ� 9{ �����8  ��������@\BBB" �������� ��������4BBBBD8 ˽������AA��L0  ��}}����lo����  ��8=??�����     `�����        ��>���>        ���Ǐ        ��>�~��>        �����                         �������         �Ù�ρ�         �Ù���         ��˛���         �������         �ß����         ??                 ���`K���        �?�����    �����������     ?�����        ��Ƿ��o�        ��������        ��������         �������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������                ?         ��������        ����3��        ��89899        ��?���?        ��������       �?8��������        ?       |��������   ""D������ݻ;   ?  `|�����ߟ�   ��������   8��������  <FBD$��ù����     !A������޾���37?ll�����    ��������s!,                 �         �        ��������        ��      ��������0@�   �Ͽ�����x  ����3���Ƅ� 9{ �����8  ��������@\BBB" �������� ��������4BBBBD8 ˽������AA��L0  ��}}����lo����  ��8=??�����     `�����        ��>���>        ���Ǐ        ��>�~��>        �����                        ��������        ��������        ��������        ��������        ��������        ��������        ??��        ��������        ��������        ��������                    ���             ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        �����?        ��������        ��������        ��������        ��������        ��������        �������        8        ?      @    <       �   ""DD          >  @|                      8          <FBD$             !A        ���37?ll            ����                        ���                                 ���                     @�      @   �x  �       D��         8          @\BBB"                  4BBBBD8         AA��L0          lo����          ���            ��������        ��������        ��������        ��������                        ��������        ��������        ��������        ��������        ��������        ��������        ??��        ��������        ��������        ��������                    ���             ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        ��������        �����?        ��������        ��������        ��������        ��������        ��������        �������        8        ?      @    <       �   ""DD          >  @|                      8          <FBD$             !A        ���37?ll            ����                        ���                                 ���                     @�      @   �x  �       D��         8          @\BBB"                  4BBBBD8         AA��L0          lo����          ���            ��������        ��������        ��������        ��������                			

		

		

		
		
				

			

		

		
		
								




			


							








			



				



				
			












			



				
							




		


										


	




	




	




	



                                	

	
	

		
	
	
	



			

	


	
	

	







		






	





		







	




	





			



					

														

					



			





	




































		
	

	
		
	

	
	
	

		

		









	







	
	






















	












	









	
	








	

	


	





	




	



	






	


	

	







		





	






		






	












	














	


	






	



	




	





	


	

	








	
	












	




	




	




	


																																

	

	
	


	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  x�8H�Z��  [�0H��B��t��M��@!�O��@!�OdM�Q�A!dQ�C!�U�3�S��S�dS�"�W��Y�� ������W�Y� �Z�Y��W���C!�U�0�+z�h@��
�
�,�
�
��
���� !�B��L��� �� ��� �B[� �� �Ԡ��!��� kܩ  [�  �9�!�:�!�;�!�<�!�=�!�>�!�?�!�@�!�A�!�B�!�C�!�D�!� � !�J	�B``��� !�B�k	�0!��		��2!��		@�2!��		 �2!��L��� �� ��� �B[� �� թ  [�9�Y[~�;�[[~�i�^[~�k�`[~�=��[~�?��[~�m��[~�o��[~�D�@W~� �l	��\~ �i	�.!�f	�%!�9�!�:�!�;�!�<�!�=�!�>�!�?�!�@�!�A�!�B�!�C�!�D�!� � !�J	�B` @ ` G g�Q�q�V�V�d�d�y�y      cb?� P(          ���  ��� !�B�9��Q�l	�1!��		��2!��		@�2!��		 �2!� �1���!�� C�� ��	�,
�	
�� ���~�!���~�C� �~�C��C�B� ΀	���L>Ü��	��	��	 ��� �B[� �� թ@P��!�~��!� �����l��� ������� �  [� ��	�!�i	�.!�f	�%!�9�!�:�!�;�!�<�!��!��!�� !�� !�=�!�>�!�?�!�@�!� �Am�	�AJ��	JJJ��	m�	��	m�	��	m�	��	m�	��	m�	��	m�	��	m�	��	� �_	�!�`	�!�^	�Z~�g	��Z~��	�C � � !�J	�B��	�5K���l	�

��ޖ	��	��	y$�� �����	����`x�8H�Z��  [�0H��B�&�
��0�+z�hX@�!Ț�ӭ%�&,Bp�,BP��J	�B� !�P�B��%�	B��� B`:�%,Bp�,BP�� � !�P�B�خ!�L1� 1�|�,Bp�,BP���� !�B�|}�<č���<�z�A�<�<ĭ�L��� �;m���9�� �!�!� �� ��� �B[� � �� �Ԡ��!�������� N�!� h���p��� ��� � �� ]� kܬ� �ܜ �� �+���4����]~ii �]~�	��\~i� ��\~� ��!��!��!� �!�=�!�>�!�?�!�@�!�A�!�B�!�C�!�D�! �� � ![�g	�,�i	�.�b	��_	��d	�#�k	�0�L	�*� �a	�	�^	��[	��f	�%� � C[���"�(�2�8�B�H�R�X�b�h�r�x� ���*�:�J�Z�j�z�%�P�B�L4ĭ�L�Ʃ��!� � 6�!�� C��~�C� �C���C��B�� �CdA��~���~L�ĭ�L�ƭN	�!�O	�!�P	�!�Q	�!�R	�!�S	�!�T	�!�U	�!�V	�!�W	�!�X	�!�Y	� !�Z	� !� ����Q~��Q~�g	��Q~�9�=�;m��?�C�F�	�m���AL�ĭ!�(� �B[� � �� �Ԡ��!��� �� k�+�  ��!��!��!� �!L~���`"� `"Y� "Ӕ"g�"��"ӗ� ���"D�~�#�%�%� �*�>	B	�
�#i �#�%) �\�� ��  �\x� � k� �K��!)? �0�0�Q � 0��I�0���0��0�	�/�"D�~�0�!�0��0�����8P������ l�l�� �� �  � �)� J	�5�j	  �"j�L8�� � j� j�8����j��!j�����  ���k�%�,Bp�,BP��J	�B� !�P�B��:�,Bp�,BP�� � !�P�B���%L4�,Bp�,BP���� !�B�|}ĭ�Lʜ �� ��� �B[� � �� �Ԡ��!������ p�!� L���p��� ��� ������� P�!� X���p��� �����L�ɩ T�!�@�(a���S ����� �,a����� �0a����� �4a����� �8a����� �<a����� �@a����� �Da����� � U�!� �(a���+a����� �,a���/a����� �0a���3a����� �4a���7a����� �8a���;a����� �<a���?a����� �@a���Ca����� �Da���Ga����� � ��+�  �9�!�:�!�;�!�<�!�=�!�>�!�?�!�@�!�A�!�B�!�C�!�D�!�E�!�F�!�G�!�H�!�K	�!�_	�!�`	�!�k	�0!�l	�1!�[	�!� ���[~��[~� C[���"�(�2�8�B�H�R�X�b�h�r�x� ���*�:�J�Z�j�z�%�P�B�L4�      0   @ޖ�V�v�v�VޖPR,Bp�,BP���� ! �ԭi �F
m 
�� ���!�|�~�!�� C���~�C�  �C��C��B� �i ��m���~�!�I�m��,Bp�,BP�� � !��� BL�˜� �B[�����p����p��� +խ�� ���!���� ���p�������� ���  [�  � � !��� B�k �#�k �i � ��V� ��"� �#�p�%� `"�� � � � H����X�~0��������� ���m	�o	�m
�o
�����
����~� �~ ���  �� � �
��� � ���?H)�o		�s	h)JJJ	=�p	�t	�
�m	�q	�w �
��n	i�r	� �i ��� ��ȷ ��:�:�	�
i�
��� e�Ȁ�� h� �0`��BW�����|z����\� I��x�x���|���x�C���������x�x~�� I���~|}��������P���{|�������� I�����~�x��|��\� J��������x�x���Z��x�x������ R���������{x�B��x�����x�xx�x� I��x��x�������x�C���z�x�x����� 8���~|����x�x�x����I���~|�����{x� @�x�������x�|�x��� =�������|�|��~�|��\� >�x����xx�x���x�Z��|��x����� B��������������`���������� ?������{������|�\� Z��������{�� 0���x�xz�|��|��~�|��\� N���~|}��������L����x����~x��� J��x�x��������x�E�����x��������|� K�������|��~�|�\� H����x���������� 8����|z�x��x�����\� C�x�x��x�x~�z��E�������x��x�x� P���z����xy|�K�x������x�x�� K�������y��x����@���~|��x�x����� L���������������[��|����x��� I����z��������x�O���|������x� I��|����|�x�xy|�E��|����x������� Q��|�|�����|�W�����x�x{x� X�����{�z|�\� C���~|�����x����� 4����|z����|���{�z|�\� F�������x�x�z�� ���������|�|�x�|x����|{�$��|�|���x�{{x{���|����� B��|��|�x�|y���� b�������� \�\�v̶����@�z͸� �$�J΄κ������ZϚϺ����FЀ�����4�rѦѾ���
�,ҐҲҭ%�,Bp�,BP��J	�B� !�P�B��:�#,Bp�,BP�� � !�P�B���%�	B��� B`,Bp�,BP���� !�B��LkԜ �� ��� �B[� � �� �Ԡ��!��� �ܬ� �ܜ� kܭ�0 ��J	)  ����@P~I���BP~ ��+� �9�!�:�!�;�!�<�!�=�!�>�!�?�!�@�!�A�!�B�!�C�!�D�!�g	�,!�h	�-!�i	�.!�j	�/!�b	�!�_	�!�^	�!�d	�#!�e	�$!�f	�%!�k	�0!�l	�1!�L	�*!�M	�+!�`	�!�a	�	!�[	�! �� � C[���"�(�2�8�B�H�R�X�b�h�r�x� ���*�:�J�Z�j�z�%�P�B�LFӜ!d�� ���j ��� ��� `� �!� C�m�C�	 �C� �C��B� `�H	) 	  ��2!�H	JJJJJ) 	@ ��2!�I	JJ	� ��2!� �!!� "���  ���p��� ��� `�H	) 	  ��2!�H	JJJJJ) 	@ ��2!�I	JJ	� ��2!� �!!� "��� ���p��� ��� `�K�� �B[����!����  �  �ty ]��  ��� +�k  @@����  @@����  @@����  @@���� � � � � � � Ā������Ā��ŀ��Ā� � � � � � � ƀ��ƀÀǀƀ�                                                    ��a��m�H
���֭ty) 
��~9���ȹ�Ս!��Յ��R������� ���(���!��`���p��� ��� �����!��b��� ��`���e״�����ؘ�-�wٜ���e�����Tۆ�h�`�ty) �J	 �!� ����R��� ���� ` � � � �� /�!� ���V���tyJJ) ��ׅ��� ` � � � � � � � � � � � � � � � � � � � ��ty) ��Eׅ��R���) ��5׍!� ���� ���=׍!� ` � � � � � � � � � � � � � � � ��ty) 
���ׅ��V��� /�!� ���� ` � � � � � � � � � � � � � ��g�8 ��  �gJ)� ���ׅ��V��� /�!� ���� `�m� ��m�g) �g�g�F�
 �ƹ�ׅ��V��� �!� ���� ` � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��m� ��m�g) �g�g
��R�6�
 ��	 ��V����ty) �'�X؅�� �!� ���B�h؅�� �!� ���B`�x؅����!� ���B��؅����!� ���B` � � � � � � � ��m�m� ��m�g) �g�g
��م��R��� �!� ����B�%م�� �!� ���B`�m�m� ��m�gi ) �g� �mgLحm� ��m�gi ) �g� �mgL� � � � � � � � � � � � � � �
       
       �ty) � e�`�g) 
��m��ِ�m�g�g� ��g���L� � � � � � � � � � � � � � � � � � � � � � � � �      �g�m�Yڐ�m�g� ��  �g�g
��R����ty) �'�)څ�� �!� ���B�+څ�� �!� ���B`�Aڅ����!� ���B�Cڅ����!� ���B`�o�o� �L�؜o�i) �i�iL��o�ty) ��Le� � � � ��q� ��k�  �q��k�  ��) ���L�` � � � À����ím) J��V���Dۅ�� /�!�� ����B���Lۅ���/�!�B`�ty) �L��Le�� �B[���� ��+� k� �����!�w ���m���{ �!�@��� � �!��� �w ���!�y �<�*n���} �!�� ��� �� �!�� ��� �� �!�� ��� �� �!�� ��� �y `��	�?���!�������L��� ���	0%H�!��	��� ��� hi  �!� ��� ���Ȁ֩  ��	:��	`���&)��!� h�	� \�!� X���p��� ��� ��`� 0�!� N���p��� ��� `� @�!�@�(a���*a����� �,a���.a����� �0a���2a����� �4a���6a����� �8a���:a����� �<a���>a����� �@a���Ba���  ��� ���Ea���Da��� � A�!�(a���*a����� �,a���.a����� �0a���2a����� �4a���6a����� �8a���:a����� �<a���>a����� �@a���Ba���  ��� ���Da���Fa��� ���8� F�!�����R ����� ������� � G�!������� ������� ���a����R��� B�!���� � C�!��� �a`� �����m	�+���o	��!�p	��!�r	���s	��� �i ��m	�ۜm	�o	`�00�-�80�.�:0�40�0�  ,00��� �:0k��00�-�80�.�:0�40�0K� @⫩  ,00��� �:0k�00�-�80�.�:0�40�0��  �,00��� 0��  � 0�0�0���  �:0�k�00�-�80�.�:0�40�0��  �,00��� 0�  � 0�0�0�����:0�&�� �.�:0� �0�0��ˠ  �:0�kh�O������#��������D�h��&�Z�� ��� �� �-"��z`"��z`Z��0� �� ����� `)���  �`)��� " ��	 "҅ ��"!� �  ��p� �Bq� ��s� ��w��  �� � �
�  �� Z� �� � `�� �`�� "��z`�� ���� 0"҅ � � �� `)���  �`)��"���` ��k�
0�� �� #�k ��Z�� i �� "���� i �� "��� `�� "��z`Z� `�� �`�� �  �� "��z`Z� `�� �`�� � �� "��z`      *      *      +*      :*      L�Z�0)� 
���� ��� `���`��� ��"��z`Z�0"��z`�>�
 �Z"��z`���Z"��z`Z�"S��z`� �����Z�( "��� ���`��`��� ��`�  ��az`Z� `�ry ���`s���e �"���
"'��"���z`��00�-�80�.�:0�40�0��L%�K����� ����d�?�f�JJ�i �  ��  
�
���I��� � �
��B �B ���� �B �� )� JJJJ(I���e)� �0 ���I��i/ e?��U���Uڊ�����J)� ���T��Sh8� )��������L}�����  ,00��� �:0kd 
 
 ��,  ��y������y�����������  ���I�ȭW���� �6�6  r㜩��y8�0���<��<⍶��L,㭖8�8⍖����w��0�p�We{�+�`���m �X���� �M������d �?�2  r�7�����r���m���� ���ζ���Z ���)� �	��$  r�  ����������  �4��4�Ȁ�� ��� �� � ��������������`ڦW�Y�W�`�K� ��k@~u� ���-�v� �������B������'��㹅� J�'�� @~�@~:�@~�'` H~*�D��K� ��k��)�����H�� � �  ��H�H�ȹ  �! � �C � �C � �C � � �! � C ��B � �
 ���Ư) ��H� H��)�0`�H�� � �  �0�`� )����� < �� �! ���! � )  �� �� �C � �C �9! ��9�L� �C �P7F� ��� C �i �C ��C � �
B �) �! �  �! ��i �C �� C ��C � �
B �i e�LQ�BJ���0�B� ��  �<	�MD	-<	�>	�D	�B� ��  �@	�MF	-@	�B	�F	�<	�5�>	�7�0`���� �UU @33�*�$  q�EU�I 8y�0�!�
=
�	{	$	��B ��P���f>����rU9�����}iVD2! ���������ui^SH=3)�����������������|vpjd^YSNIC>940+&" ������������������������������������������}zxvtrpnljhfdb`^\ZXWUSQPNLJIGFDBA?><;9865320/.,+)('%$#! 
	 � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �    � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ~ y s m h b \ V P J D > 8 2 , &        ������������������������������������������|�w�r�m�h�c�^�Y�T�O�K�G�B�>�:�6�2�/�+�(�$�!����������	��������� � � � � ���������	����������!�$�(�+�/�2�6�:�>�B�G�K�O�T�Y�^�c�h�m�r�w�|�������������������������������������������       & , 2 8 > D J P V \ b h m s y ~ � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �      � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ~ y s m h b \ V P J D > 8 2 , &      �_ 0�PX� H"�/H$v	H$H$i �j��#W�"M�n�l�l�<$KH H�H  H �H � H � � �H >H ��H$ H$� H' ���"�#H �P $V�  �Pb<3�A$iA$vA$�A$	A �A �A �� Hr$H�sx X�{��_ 0�`Y�   � � � � � � � �Hp 	Hz Hp Hp�Gq�oGx�!�p t���t��t���t��t��u� u���uf uV��uW uY��uj u���u��u���u��v��vg��vh vo� v��v� v�� v���v��v� �v��w�� x���x� x�� y���x��y� y���y��y� Hz�Hz,�z s��s� s���qU�hq]  �q7hr��re�sUht9 hu �u]�v'��v)�wH�wV� w�P x�Phxh hxm hyc   r���r� r��Hr�Hw�hs}   s�Phss  �rPhrt  hq~   zrP zvPAp�Ar�Aw�Az��p
(zK$��l�Ppy �Pp�Pw�`��P��P��p�p�p*��p��p
�p��p��p�q�q	�q�q2�q2�q�p*�q!�qB �qq �qr�q��qW��q��qX�q��q^�qv P�o p�o qp� `� �  ]t� ^� �� ~� O� O�E� ��P  po� �� �� ��0�!p�!��!p�!|�!��!�	�!��!��1�1&�1F�1g�0
�0�0� !� !� ,� �� 2	� � � � �0d�0d�1`�0��0u
 !�p�!�	�!��!�	�1��1	�0 �0 �0,�0\�0� 1�!� �3�3�3��3�3"	�PIp�x
q�) �-)x8 0x	 !�x1x3: 3x6 �\� P(@ � � �H  D BEwH  �w�H @H �H � H�H �C $H(C)� %N� H�Hh Ny HO H� N� N� H� H�H�H�F� ������F� H�	H�HjS ���H"C,�-C%H&C(�)C%i&H& C,�-C!�d�j�Z
h� h� H  /H  	� ��"�H".	H"� l!& l!� H � H �/� ��"�Ht Hp AHp 	Hp�	Hq� Hp�Hr�	�p��p� r��Hs��s�Fs��s� Es}Ds�Hs�Hs� Ft�	 Hs�FTx �Tx�T��ET[HT HT HT( HTPHT.*Hc�T���HT�ST��TR �T� �dM �d� �d� �td �tE  c��Ss��T���d��tJ��� t��Ap�Ap�Aq�Ar�	As�As�As�As�At�AT�A �A �A"�A �A�A�A�A�A�A�	A�	A��T+  �T�id)iTlL lE Hd( Hd) hdU  �x y xp"x px+T�J �����`  � � �!`)A�!e&"i&"j)1k1l2cXA� 1Q1�A	A�g1� W1�WAWAqWA�c1�c1�c1�cA(cAV1�2�1�g1� gBp W1�W2�WAWA<WBAc2�c2�c2�cB$cBGcBucB�2I2�2�BB�BZW2zW2�W2�WB,WBlBYWB�g2^ W2�WABcAy�1���A*��2��B(��B� W1�!�!�"�X1 !��B�8 ��_ 0�PX @F0 D1%E1.D0&�0y��0q�2x��D2)�2xH0 /H0 H0pA0�H0�	A2�	H2�H2.	�0H1�A0�A1tD0�H0� H1� H0�H1� D1�H1� H1� H1�A1�D1�H1� H2� H1�S0�S1�S1�S1[H1(H1JI07I2:I1RI1_�2�M �^�J�p`�d H@ HA	HP� ���_ 0� X��Hr*
Hp�/�p��r&�rWDq_Dr'Drx�q��p&DpG�p���Hp� Hp�Hpl Sp�Hp\ HpO Hq~	 Hq�	 SrFSq�SpS p�2Pp� p�5Qp�Rqg� q�7Qqh rh4PrX  rH2 q�4 q�2 q�:Pq� Hp 
Hp /�r��r��r��r��q#�q3 pH? pY@ qr? p�< q�C q�D p�? q�A q�B q�E q�? r7?�p#�OBe42e44e461&�������� �"��J��8�6��?��D���O�e���l�������:��&e�e�e�6e�8e�:��#��e�1�rOJeReR�S�S�S�S���������b�v3�n�v:ak8��49S^p�X�F�=�e �j���&��
TT&&G��/&�5�I��;¤Ke�Ce�Fe�Lk��D��M��>�P�L�� � z |  � �' r+1�-��tچ!ڎ+e|e�e|'e�%Of��rt+�l�z�z�z!�hjnjnjnOj��4�H�����
r�r�%�%���#��!��%��'����(D���,������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������1�����������01YI           YOSHI'S ISLAND         3 ��,O�O�O�O�O�O�O�O�O�O�O�O� �O�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 H�����0       @ x � � �          � @� �               @                                                                                                                                                                                                            x H                0          8 l D               8                                           &                                                                                                                                              �? �� � � � � �                ��������                                                                                                                                                                                                                                                       #                          0 �0�                                        � � � Հ׀�����@ 0@8@8 ( (   �@�@������������ 8   > 
       ` � � ����׀         ` p p (_ > >.&�@C�� >                     �p�                                                           0 �0                                                                                                                                                                                                   �? � � � � g             � � �� � � � � �              @ � �o�m�#�#@    0         �����@�������p� | 0        � ��������v���              �ց��ԃԃ����� � ( x ( ( 0     ? � ����@?@?@?           � �� ������ � �           #�?@�`� � ��g�             |�� � � ���`             @ �  ` �`��d�| �           �                                                                                                                                                                   � h             o               	 �   � � �       L0�|� � � � � �          0 �     �p� � ~ <�{�1� p     � �    � B�<��( ��<~ <    � �   �p� � � ���� p         � � � � � � � �                 � � � � � � � �                C Q ) &�"���� � � � A A a    � � � { 3   �        � � � � 7 � � � � � �               p � �                                                                                                                                                                                                                                 �          � �               , �        � � � �        (�    �        � � � � � � � �                 � � � � � � � �                 � � � � � � � �                ��������   0 0 0    4             �q� � � ��� � p                                                                                                                                                                                                                                                                                                                                                                               @@`/`/p?    0 0     � � � � � � � �            ����� � �@�               0��30� � � � �                ���`d��	� � � �                                                                                                                                                                                                                                                                                                                                             < �< � �                p3p0p0�`�`�``��         �               � � � � � � � @�@            9�?��� � � �  { 1    � q     � � � � �� �  ��  �g   � � `� � �                                                                   3                        � � ����                                                        � �              �                                            � �              �                              @@?�?  9�        @ � �   � � � � � �`��o                ����� � � �                 � � @ � � � � �   ?�                � � � � � � � �                 � � � � � � � � � �� �����                                                                ??g>�~>?                ���������������@                  "gz      ? ? D���}	����FS�x � � � � � � � 
� 0��         "��A���r��#�< | � � � � ?    	�����       ���F�� � � � � �             0 ���� � � � ~ <            � � ��? ����              � �@    � �����?��@@`                   � � � � � � � �                 � � � � � � � �    @@@@�����0� � �  `          � � ��                     88|8|0                =;�{���o                �`�������������                ?  	  &_ |       0(  �$� �?� � � ��~� �  �       ��� ����[�  � � �    � ��m � �� �D�� � � � � � � � � � ��G �`� � �������    � �� � � � � �               ,�? � � � � � � �         �? � � � � � � �              ��������000                � � � � � � � �            � � � � � � � � ���? ? ? ? ? ? ` ` @ � � � � ������ p p �p�p��                �t���h|>>O>�                3s????�;                ����������������                |x�	xt����03 ??    0<C�� �`�@���?�7@À�@���@� `00 8�~t�?����>�~�  ?  8888@�G��@�@����~�|�� �   `�����/`�p�p����0 0 ������ � � � � � � � �           � � � � � � � �                 � � � � � � � �         ? �������l �                 � � � � � � � �    � ��� � � � �  ?    ������ � � � � �  c  ~���� P Q                    >>���������                �{;��ߎ����;                ������� � ��Á                ��������y�w��� <? ?   <�8�G��t��p�8�0 ?��@��@� x 809�]�]�+�k�w�o�W�;\\\\((hhpp``PP88����������������      p�p��`�`�`�`�`�`����                     � � � � � � � �             � � � � � � � �   �               � � � � � � � � � � � � � � �                 � � � � � � � � � � � � � � � � ��               � � � � � � �                        ����?�?����~ T              ���������_��_                � � �����@��@�                 �xtxtyw{< ??   �00�O���@���� 0�� ��� �   �7�;�;�?����00 � � � � � ���������������@         A@�`�G�>� � ���  ? � �   � �o �	� ���@�� � � � � � � � � �!� �� ��@�� � � � � � � �     � `�0�8�x�� � � ? � � � � � � � � � � � � �     0` �@��� � � � �  ? ? �0 0          x � � � � � � �   � @   0 �  � � � � � � � � � ����������                TT�@�@����x���            �?�?�����?��                ����������������                7	         �?�? � �@��3�� � � � � � � � �7�7��O��<��  � � � � � � � ����ǀ�       �� � ��.�-�3�3� ? ���Ȯ�--�����@�� � ��ýǻ��� � �  ����������� ��s�j�Y½� � � �ssjjYY��� � � � �@8�8�8��g`' WP������  � � � � � � � � ���� �� � �{ { � �  � � �    � �� � � � � �  �     � y���� � � � { � � � ����� @�@�            ����      ����@�@            @@@@        �������?? 


          ���������                    (x�?�q� ??������� �>� � �`�   ����������� �@�` ��� ��3 �@_``����������� � G�G�g�w�?���������������=�=����6�u�s��==���旗��uuss���������+��������������##������½ü���R�����ν�������RR������8�8�� �����=����  �� ? ����� a���w��     � � � �  � � � ��|�z�t�h� � � � | y s g  � � ��?0��� � � ? � ' 3 �  � � � � � � � �� � � � � � � �                                                                                                                       ��� �w    ��������  l����� �� ?��������������??�!��� �� � �������������������� � � �    ������������    ����--    ������==    �����<��[�mm  ����<<��[[��  �����{���]����  �̳�{{��__����  � � e�e�=>  ��XX����   � � )��/�?�6��@  ����&� � 2>a``p<   > ? ? ? ?  '&;>������� � � ? � � � � �  �  � � � P��� �         @� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     � � � � ��� � �������	�� � � ��������
�
������ ���������
������������������������ ��
���!���
�
�!�"��
�
�#�$�
�
�
�
�
��
�
�
�
��
�
�
�
�
�
�
�
�
�
�
�
�%�
�
�
�
�
�
�
�
�&�'�(�
�
�)�*�+�
�,�
�
�
�&�'�(�-�.�/�
�0�1�2�3�
�4�5�6�7�-�.�/�8�9�:�;�<�=�>�?�@�A�B�C�D�8�9�:�E�F�G�H�I�J�G�K�L�M�N�O�P�Q�R�S�T�U�V�W�S�T�U�V�W�X�S�Y�8�9�:�;�<�8�8�8�8�8�=�>�?�8�@�8�A�B�C�D�E�8�F�G�H�I�J�K�L�M�N�8�O�P�Q�R�S�T�U�E�V�W�X�Y�Z�[�\�]�^�Q�Q�Q�R�S�E�_�Q�`�a�b�Q�Q�c�d�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 ��   T         P                     U   �       �Q   ����������@ &XP   �      n 0                 X                  �����           ]~   ]�             ,�Z~��~�Z�             Z~��~Z�           &�\~ ~�\�           &[~Z~[�           �[~�V~�[��          \~�Q~\��       �yw�M�2H   B�        �  �                      � � ��1                  <  )�#�uқ�����  �� 8    �   �  �� �  �  ( (q q  ((                                                                              �                             1                                                                                                                                                                                                                 _� ��w�                                                `��0�0���0�*�������� � ===���=  OҦѪє���      ՟��ԧէ�     z Q 4   Q z                                                                 � H�       �                                                                        � � � � � � �`w  � � �       L �9�Z�Z�Z   x   
    
                    
    
    0 ( 2 0 ' 0          � n�            < '           $�;                                `�                                             @             �Ͻ� ]������ � =��� =���?�
�H�`�?��?��<�]?����� ��� �S��� �
���iML��L��� �']��� ���E�F�D\\�kk�� ��m�8�`�C�C�#?��?��?�?7!?f iML�����\��L�S��`�Q�Q����?T� ?�_D��� �G�1�?F==G��_D��� �� u� ���� o��� �� u� ������� � o�ʐ?����Ȱ��$G���(`�P`���a���`��\� |ՠ� ԰� ����	G^	GE��Ԡ���ԡ���
�a����a��`�a??5� ���4�	�����z�M�� ��]�3��2��5-�4���ݍ z�+�/K|=������ ���� ��m�!��z��!����z�}�\��?���-�G$���� �� o� �,?��<?����\?�?W� ���� � � ��֟��ox��@�Z��� �[��Y?@�\_[����Y���p�Y_[������Y� ��_[oh���h��h���h���h��#h��h��	h��3h�Qo���S� T_[��T�D���T��U��S�T?@�V_[���_g�H�F � � G��Y� So� �@:@-�@:@��o`� �����]������o����@��H�F o���G�G$(��#����
?
	�Ձ��Հ������Ա��KG���Z�h�T�P�B�_��Y� So� �_p������_���Yn�?����_��B�B?��B���@/�����0 ��� �G�1�
��� ?�� Ԁ-�G$(���ԑԐ��p==G��� �^�G�D�1�n�p�d?����?+
�����0�0�1�1/�0 � ?�0-�(���?��(���?�?�h��?�/�-�G$��?� �p�������q/?g?�
==G�_��T��VzRnT�T�R�h��dz`�`�fzbnh�h�`�j�b�Z��\zXnZ�Z�X��^� �G�1�?�==G��o���
-��
-�\��2��0�0��1�o�����`�_���`� �=�$G�:M}�\]� �(8 HH 	GI�/�GNI ��� �� =�������!��� o�Q(�1� �0oԑ-?��P��1�?@�@��Aoհ?�ա?�Ա��� ձoձ-� ��Ξ�D��o���	���� �Xo�Z?��[��Y�Z?@�\o� �R��o�T?��U��S�T?@�Vo�Po���������o��?���?���o�/� Ր�Ձ?���-�G$��� Հ?�ՑoՀ��o�� � oԐ-?�� ���?@���o�������Ձo�@?��A?�Ԁ�0�0�1�1�@�0�A�1o���J?�� �`?�� �b�Ho�h?��i��a�h?@�d?��j��c�h?@�fo�`�b�Ho?�
?��N?���]���?�=�`����Do�M�}�� �� dM�+(H��L`�L�L���� � �� ���H �l?��M�}?�H���<�m_��_o-�G$��&�/���D�0h��>�G$��?�n�/-?�?�ԡ?�Ԡ?�`�P��(Հ��a��m�?@�p��qo�a��`�o�kH��� �-� ���D����o�
		1	=	X	g	y	�	�	�	�	�	�	�	
H	�	�	�	
6
m
t
L
�
�
    ���	� ���?C���#����	G^�����/`����?�/����?����	�0���?C�G$^�I�1��0�}�\�����������`����P�!��QݐH���?��� ���3�o	G^��M�`�
�� ��/	�?`����o�q�e�q���p\���0�1�� ��0�0@��h��?h��)h��0m����
�/���#��
�1-�0�/��A-�@�/���-����/��G�\?����������/�$G���`���?F?5���L��ްD� u����/@�  ����`��Ա��`��ՠ��H����h�(�/�ݍ ?�_o����o����	����?��1��0����
�A��@?��?�?5������
�q��p?������ް��Q����`��_"��?Rm�Q��� �Q��z?Rz�o��Q����`���H�����H��Y���������!o )4BQ^gnswz|}~       X����!++���43 ����,<MlL\=-\acNJHEIKF_�e	�	�
,��J���*Ver S1.20*��� ��� �� h���/ �� ��^� ��� �� ����/��^� ��� �� ��� �� �� ���1�� o             oohXmhXMLXXXXXXXXXYHhXnXXXQXhhWn////XQN////////^nXXXXYhhWXXh^hXhXXh?hhHHh>hhhhhhhhhhhhOOEEUUUUUUUUUYUYXWWXXXXHAn?nmnXXX^^^]^^?????_^^^^^^^]]]^nn^^>?NXnE^XnXXXNHXX C65I56-N??O_F5mF^N>N9MFF?Ihh^nF^NgLE9MFF��d�&��	���������=dz���*:����ctc:F�SY_ekqw}�������}n�����CI"9cY�z)e5hmIS]gq{)3!��7���������K�������  ���t�YaSx(�Rd,\��������z�e��@8�LT�a6e�Zixx���    c          I        ��cc���H�*/IWfu�M���Pj5)/IWf�d�� �Y� �d�� �Y� � �P�� �	Y� �F�� �	Y� �<�� �	Y� � �o�� �w� � �d�� 
��� 
��� �F�� �(�� � �Y��������M����F����?����8���� �8�� �8���� �	x���� �x���������� �x� �	���#�#�*� �Y�����$� �PZ��
�� �F������������������������������ �d ���� �P(���� �<<���� �(P���� � d���� �d �P�F(�<2�2<�(F�P� d�  ��2��(���0 � �P��<�� �Y���
� �Y�� �Y�� �Y�� �Y�� �Y�� �Y�� �Y�� �P�� � �F�� � �<�� � �<�� � �F�� � �P�� � �T�� �� �?� �1� �#� �� � �T�� � ��Y�� � �*�� �� �1�� �� �?�� �	� � �T�� �� �?� �1� � � T�� �� �?� 	� �F�� � �t�� �� � �T����F��8��*��
��
���� �8�� �� �48� 0� �d�� ��� � �� �� �	Z� �Z� �
x��
���
���� �x������������ �	O�� ��r�� � �>>��E7��7E��L0��0L��S)��)S��Z"�� �x��z��z��z� �T�� � �d���P�(�� �	x�x��(� �	x�� �	x�� ��x�0x� �n�� � �x������������	��� �x� �x�� � �x� �x�� � �
d�� � �d�� � �
2�� �2� � �x�� � �0d<�� 0�0PP� 0�0<d� .� � 0P�� 0�0d� 0�0x� .� � 0P�� 0�0d� 0�0x� .� �`P�� `�`d� `�`d� `�`x� ^� �`x�� ]� �`Z�� ]� �`x�� `�`� ]� �$x�� $�`� ]� �$x�� $�`� ]� � T��F8�8T��*����*��0� �x�� ��`d�� `�`� ^� �0x� �2� �d�� 
� �d�� 
��� 
� �d�� 
��� 
� �d�� 
� �d�� 
� �d�� � �d�� 
� �
d��� �Hd� � �H
(� �x�� �� ��� �� ��� �0� .� � �(P�� �� ��� �� ��� �0� .� �0n<�� 0�H� H�Z� X� � �0<P�� 0�H� H�Z� X� �<�� $�$d� $�0� .� �d�� �� � �d�� � �d�� �� �d�� �� � �d�� �� � � �
(�� �� � �d�� �� �d�� �� �d�� �� � �2� �2�� �x�� � �x�� 	� �d�P� �d�P��� �d���� �F�0��*�8�?�F�T�Y�T�$�����0� �0P� �T�� �� �?� 	� �0P� �0P� �0x� �0x� �0x� �0P� �Hx� �x� �P� �P�� 
� �P����� � �P�� �� �<�� �� �(�� �� ��� �� � �x�� ��� � �x�� � �x�� �� � �d�� �� �d�� �� �d�� �0� .� �0d� �d��� �d���P�<�(��
� �d�� �� �d�� �� �d�� �� � �x�� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� ��� �� � �Z�� � �x�� �� �� � �x�� �$� "� �x�� �� � �P������ �0P� �P�� � �0x� �0x� �0x� �0x� �0x� �0x� �0x� �0x� �$x� �x� �x� �x�� � �x�� 
��� 
� �x��� �<�� ��� � �x����d����P����<����(���� �x����d����x����d���� �x��� �d��� �x��������Z�F�(� �x��x�����Z�F�(�   ��x��(�  ��x��(�  ��x��(�  ��x��(� �Z����d����x����d�$(� � �Z����d����x����d�$(� �x��������d����<�$(� �P�� �P�� �P�� � L��7��)��& ��L ��7"��3)�� 0�� L��"7��3)��0 �� d�� �� ��$d��������`�� `�0� .� �$d��������`�� `�0� .� �$d��������`�� `�0� .� �d�������`� �d�������`� �d�������`� � K�-�<� K�-�<��$d��$��`� � �<�-�K �<�-�K ��$Z��$��`� � �-�8<�-�<��$Z��$��`� �p �8 ��$F��$��`� �n� �n� �x��� �x������� �x���d���P���F��� �x� �x� �<�0� � �<�0� ����
� �� ����� �j� �j� �j� �j� �  jp 
��pt�
�p �jp ������p�����0 ��������������@�� 
�@�t�� �� �� ��� �׸ 
�Jp 
��p 耍\?���(���J�M?�� ���?�� ����ĮĞ��ŏ��Ŏo�@؞��� �.����?@�����h�� ����?F��/�
�_�� �?o���� �	~����	��� D(�����-/C�����
/������Jo��耍\?��� ŎĮŏon��?��?y>�J�J�M?����0Į� ��(]� ����D?o���&�?_>���/��
�_�?��1��0��?o�� Į� ���������pĮ� ��(���D?o�(�`<<<<]��]�t���?�=�n����/=���.o	  �   � p   ��	  �    ��  ��
  �@	   �����������������������(����]���d��_�>�֠��K�n��������_� �� e� ���� ���.� ���h��Po� Ű�š��ı�����  o� Ű� š� ı�����  o���� ��?�>/�(�H����\?��/_$ ?�>���h��h��ՠhp�hr����  /h!�?� h"�?� �ա� ՀԠՁ���� � ���\?���]��>�Пo� ���,��@�������}�\��������_"L��o�����ա�_d!�����~Ց�-�}Ր�,_8"�~Ց�-�}Ր�,_8"����hp�	hr����  � ՠԠ������Ձ��Հ������ ���� �D�?���%��$J��J`���J�M?����������o?�!_d!?�>��������,���հ�_�":,���\��� �,��06��ֱ:,�,�0(��?�� :,�,]����?�}/���?�� :,�,h��_ >h��Gh��X���?��?y>����հ������?_>/�u�����\?����-Ց�,Ր_d!� :,�,���D�?��?y>� :,�,��ԡ� :,�,��Ԡ-� :,�,����D?_�"                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              b&R&  r&�&�&�&�&      '              ���������}���|���{���z���y��F� ������}���|���{���z��F���$����}���|���{�����F���6����}���|��F���H����}��F������������
�   '  0'�'�'&(        �����`d���������� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� � ���������� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ������������ ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� ����������� ��� ��� ��� ��� ��� ��� ��� ��� ��� ��� �� ~(  �(�(�(          ��������������7��{�)�?�9��� �������������
������ �(  �(B)�)�)*>*y*�*�������	��2S�.w�Z�z�4�d�6�5�
H�F�7�h��I�(�)�*�z����* ����$�<Z�C�k��V�8�
Y�6�S�5�
X��g�i�I�9�!:�0�0y�F����	���T�J��;Z�z�T�4�Y�u�V�x��
V�x�	�9�7�:�*�.�t�.�������
���Z�8�0�*[�z��i��	6�8�	W�V�	Y�v�Yȟ9�Z�%<�.�t�.�������	���o��.m�e�x��d�J�L��{�`����*����2�.��i�l��|�9h��
j�
d�
Z�z�	Z���
W�z�-���*�����w�z��/{�w�I�J�L�{�Ei�	Y�
Z�z�i��V�v�`�-�3���
���b�K�W�	R�-���%B�`�.�2r�+�5� ��������                                                                                                                                                                                                                                                                                         X�n�P��n�	��
\	�
�NP�� 8 ��8����L�\�
�������J�<�H���p�8��\���l��j�R��n������F�����&����������t���\�������t 4�b�~� J2��tH ������� ���� ��������"���@���(�����z�<���&�� �$�X������t�B ��.~
j��tLhH�`	�������X��4	��������*f����t�������z���f�l�����t��z�^������6��h���h�*����������:�*����n�@��� d�� < `
fF���8���Z���^�����������(�D���j���\�������p�������l�������V ����4�� ��r���D��T�"z��F�����b����(�����������x�������4�\���� ���,�����D�,�V��\���l�`����F��L�����(�F�z���H�F������T ���F H�f � ��� 2�v��*�����Z���6�8�l�V������������������V�����2������d�������(���P����� ��������n���<���������l�f� @���:�������0���6�����jPdr����^J����	�����>
�>j��n �� �n
��

 
���2r�D0\���� ��8D��N�&@�,������>���N���b���F��<�~�V���:��z�Z�����f�F�����p��D���B��$�x��v����8 P�  �D�
���	����rZ
����H�����	���tj��������h ���4�~$����$ ���������$ &�� H�������X�v�6�����|������
�������V���f�����~��n�z ����N��� ��������v�,�*����~ �Z d�������
� D��.	��
n����\��4�>"@|$|�vp`D*`,.<T��� ���
6��	L�>z��
J����\���������z����
�r����v�F�,���r���Z����V��� ��\��� ��>@ �
�
V�	60z�*>0��N��v ��
� ���~���.���b���f��XN
<
���&Z
��Z>��lP�&�z	���* �Z����nj����� �������R��l�����N�|�h������� &�&��	�nN��z��R�.���~DX��"������b�	�
��������d��p�X	$��v�������� ����������$�h���X���,�J������&�&�p���R ���\�@���@�~���������6��, \���j�r�������*�� ������� B�����"�.��� �B���� *tB�� �� ��|��F�B��F��v^:���&�
�&
&� V���|�����j���\� �(�����J��2�v�`�b�H���b�z����������B�t�����X����*$�^D	�r���.���R
�R> 8��zrn�� ������F ���B�t���r�~���������� �j�2�������������������B����f�� ���l���P�&�0���������f������H��`� ��������������������$���<���j���T�@����>�����V�����t *X�d���B
��H

���
.H8X�X��������4��xt����P�~ ����N~�@� ��&�>� l�*j�� ��t���~������B���4���v���$�n� �����F�������`� *�v	�8	���v����� ���h�����t�P�4����������� � F�����4v�Tn��� �R�	��	� ������������*�x���� 8����� ��@���:�������R�����������8��"�<��H������V������������������(��� �,�f���\������   P�� � ��� hN�N� Z��������@�����R���T�����.�H���b�<�������4�
���2����b���8�����������f�P�D���� <�* �� �.�����.���|���"�&������~��� ��������� ��N��JB
v�V`6�	��^ ��������p�� ��t���������� |B�r�Nz��J�n &(� ,��`�z��<��4�,�$�����t���@�L�J���������\�������v�f�����N�f���������b�p������ �T� �� � ���
V������|^N
����*p�p������@R���l�T�4�f�r������ ���|���"d�����x��r�V��R ����H�� �d�H������f� �\�8���������:�X�"�������L�R��������d�&���������@�f~�.�	�������z��	�,
V�Z2	J
,LVN��P<P���&l�z
�Z
��	��HrN |������� �����
�����*�L���>����������\�F�������B�n�z�P�������F���Tp ���&Rf�����8
��
�	� �r �r �� ��	� p
� �	��	��n
������	���!rv#��"Rd"�D!&�LFv�����$�N����TN nz�� ��$���b�� ��P�4���������H�Z���@��	V�HD��� <h��>0�nJ�z� ��\�d��x 0��hB�HZ����
p��v���h�����j���,�D 4��V�������r�:��:��
(|	���X� D4�� J ���h<���@ ����p����"������<�f�|������< �H � ��X�H���v�:�2�����L ��� .�V&�6 �� �� � :�Z��	�H	jf
�*���
>$d�&��:� ������R�����������*�����$�X� ��������V�����D�^�B� ������V�|	DlN��� X�	��:�`������������ �r�D�Z�0�������8���`�4�6�J�����$���"�H�B�Z���������*�d�4��� �������@����� ������F�|�������d�,����,�����������p�2������2��^�����"��������h�N���`�Z����V������R���R��L�	2	`l	V @@�CGYGY�d�dIfmf�g�gllgl�lWpWpMwxxWy�|e�����8�8�����z�����������ʢ�V����䩹���u�u���`������)��                                                                                                                                                 ���������������
����� �����
	���
��t����������� ����� ����� �����z��Z��?�������� �� ��=                                                                                                                        � :,�,�Ϗ�ҏ�z��ҍ ��]���mM�?�m��=�n������!���� _6"��`���?F�a��`�� G_o-�\� ?���L_�����Y����Yo���
���Y� ��o��$J��J����J�M?�o��                             �      �          �              �  �                                 ��     �  �   �            H}       �    � ��  � � �� ���                   ��    �� 0        �  � �                                                                                                    3f�����3Lfr����������        ��2�;�<�.���,�>��в������"D�S�Aİ9�β�$�Q���"� E���� �^�_�/�Rв/ �a3��o��������@��?��/��-�V��3��. ��]���/�]�L�?����.���_���o�O��� �_O2Ҳ*��00�/� �D#�6SC@u�������11���.�����>�_�A��B �#<����!�B�?���#����R�!�����/$�/��ܭ����̲!!��1�-�CP��,�'+������ ����2���/�#"P�%��!�5��`� �-��"��4�=��#-������$�T��F�-������ #0����E�>���˾C��������� ͢��O�2/� � ��A"<����S��!�T���O�4=�RS��#���ܲ� #��P�?���. �   �������� N���>��!�./��M���=L�N � ���жm��f�� �[ ���1%�!�����,?@ ��������m��!�M�Q�  Ϣ@O"�,���� ��"���4� �3�������4 �]_#=��\��Bղ��2�l���N� ���-����!!%�������-������M�1"�SVCJ
�/��M�C$����B�O0���0�C���.02�d$� P��!���J[�����" ���M�@� �@�K��=�$��϶� =M�]��`��:�������!�M#���?���p����@��" �OB�����1� �"��,TA���R��0�������2�;�<�.         �O-.>>/t�c>���x@�"��.� \>���AO0��� 22�����bA�ޔ��$"������U0 �̘!-?]�����db �����ߔ��TR!ڔ�� �ϔ�Sr?ڔ�"#ꡨ��N<=�m} ����PP?�N>�PP>��!" ���Q`/��#%4/ɭ�3C�� �����.#4̤��� �ΤDB ܘA!����ԤCC ܤ��Ͽ� 5C �ۘQ}2ᡣ��.UB��ܤ�!#�͠� _+��2!2/��¨��m�� 21"/�˳���]� �A����E��V���Ϥ#B"���B������#2!켢Q�B ����E!�����>�#��A�BT�#�� ���! ���@/�2�� ����  �] "��?� ���A �U��/��&!�����OS�]���$e���$��3�ܽ��EP����@S>����2A�����P%0ޤ�,��W�-���$��B����3/��� k  ��_ ?���OU>��� Q�����L $�����#��2�� ��3 ��� ��-��/��!����]�!�^�1�O6�n��+�5Q� ��O��ߤ��-��D�� ����C����"����� c����e!�1ʸ ^�"���2!�ݴ�^ U.����4B A
�۴Q�&0��.ͤ3#��G�������"���.�.�/�����N�?�? � ��>d�=� �# �!��oFN���! ���P�6@ޤ���E ��\�4�����ܴ�P�60�������P50��޴�" ��P�3���"���P�4��#Ѵ��OD�m���%4� ��NU>� /1 � ����Nc���1!��>����bB!.�۴��S�� ʹ�1!��2��������"��B����� ����L"�^����$"����/_ܤ����T3 ����d���\.���A���������P &O��ߴ���>�0^�  �@N�������.���m�$���2�%�����OV=�Q�B`����-���$N�����]����"���N�0^�? � @�" ����c�� ��2���[2��3�C����7�N����T3����m�����!/���0^�!� �3"���4Ѹ���-��/���^ e�,���#�� ��5��Q͸������oU,���$� �δ5��R��ϴ1/���^�u�� #�����n����"� �F�=Τ�!��TQ�޴��oU,��
�F��˜�o��΢!-��2/��� �L�"�?�1����N e��!�?!�и��y�4�����%ͼ��U�@��.���-F��r��� �A ����>�}�2 �/O������}U�3C�]Cѿ���O #���N�����@ �������A����!������B��� ������2�/� ��c��ڭ�A�.�� �!����A���������Q��� �����@��.����O #� �����O �Q���C�����^ c��4/�����1���� ^�/V��_� ��!��A��;�  ��2�����o #��/"�����/B�� �3����%)�@?��L���Q�#�����V?����/1����2��4��/� ���# ��%��0�!�����1���c,���C�.� !���!���^ �3��/�#�� ��0Ͱ���4O����`�$�/������/�.�0�N�� �B�.���%�E-���O3���1��/�D���0� #������1��?����۲!E.�%�S���"R����3���  �N�A�� O����b�.ϰ�5�U����N2��.�1������@�.�/���1%Q���c�S������U���"��1�@�"�2�����f�*�>�E=����1%P��B��1�������@�#��2���B&�_��A��1�� �E��/���2������ O�B�� �/���#�-�0������2V���!M���1%P�1���1������P ������ 6Nߴ:�U�A��"R��"���2����!�A��1�����A%N��4=�&�"��� �e��$��3���0�_�S �!?�����Rݰ�V��d����! E-�/��&>��b�3�!�������e��C3��P����Q$=�0��"���C��C��#�3����!�E,�$2�S��0��$�S��$��2��� � 4-�0��/���S���U��cٿ���"�U,�#�/�� ���E��3��2���2E�M�/� ������E��]�6
�U߱�2/2��2���!����"��4,� �#.����!�E�q�O���B.$P��1��1� ��2��E=�#/��/����D���U�T
���B-a���!��!����2DN��1��1����"��E-�# �������5-��5N�5=����E����"���#� �C��"��"���B.�A��"��"����R-Qް�D��Cھ���AQ��2���!����B�A,���!����A�,�������R.Rް�B�C����C/�C��"��2� �3� �C��!��"�����E��" �"�����F.�Q�R��@���3�4=��"�����14N��"�����A.�2-� ����C/�D���S.�3�����5�C�#/�����"�D=�������A�2-�����D���"�0�� ��� ��24N��5��#�����B.�T��.��/������E�!������1��4M�����1�S��!�"������5=�c��#���"/�C��>��B��1���!�4O�������3�/�U��2��� ��2��$_�!������!�E���B�1���NAѰ�0�������5>����# ���C�!�!���!��������!�!0��������E��!�����c=�C�    ����3/C���A� ����# D��M�� � ���!C��L���>��" D������A,��2�>�AѴ ����_2-� ������"� �E�� �������4����@ �� ��N�a*� ���C��� 0� �  ���2�d:�����ٶT�>�`?�0�3���A�2����Eo�C��������2.�/�� ������en�D����� �f�5n��"������T��3��P��0�����ܳ�2?����5=�����6��1���@������"�F@��D�0�̿���<�#Z�C����7��E��-�!����#0��� x�nm0Z���"����L��%�@� �"x#$�a�x���P,3t��@��t �D+�3��dFaOˮ �Rt1��<Fp$3����d��12�h2�A���t!N ���`�#@,��"@hL���`h?�����O d3.��/�Cd��%p����A��`.�50U��hJ���J!�d��O ��d@,���#�dN��?��dB �>T.�n=�T��-?��$T�2��U�"T*�f��A�d��st�dT������0d�+�4!!h���-!�x�A �����������ё���%��!�Ӕ��0"!!��������ߡ���P�L=?,�N��QQ!C0ﭘ�l;>\+���߯�%�������������/�O> ��4�������� .A�!�:_>?�0�?-K.].%�2���On<.�!� �FS?>=�)���DrA�2���!3�\��_�Ӕа�$"����R����ܘ0�B�"O�����τ.�=@6&����A-�2 ��=�?O@O-��lA0������Ք6����;ʤ -.1O�1��0��P.@�-1�����A.�""������NK�_1 
-����%���ޔ�</A3� 
����ӄ5c"̡ބ��""F3������>�4#��Ҿ��"/11�>��Ѳ��Ua\=����B Q/�/���޲-�#R<0������������"��=,�A>"���\}]\�)�M*�1�? BN. �����Dx�0>��OY�4��E����������1����!M�� ?LNA-�0??-�����a#^�ΰ�D@��"�m�=��1C���ñ����4�4!�������B�+�������T��1�����t�"S A���Т���1�N/A1��݄����t������	ʄ -�C? @x> lZMx?!� K t��۽���x䤷���\jt�����ń���h�][�.LxK.!���x1����d�m� �x<[,O?�#�x�ߴ�-xM>��䳴�x��6��QhR���_tN/!�x�//-?xO �x� �- h�󥥦��Qt0�����h�š�_�6x=�����t !A2.�!t��"�����d���$%0�Bt�����d��a?"D"t�!���t������d�M".�/d���-!Qt� ���d㞰.
�Dt�3?�$.�!t.�./dR>3��dA�1<���t������h����@�d��Q=T-�`&V��#��t ���hD>�T���d ���MT$" B*dN,-N,/T��0�6�p"" ���Ͱt����.�e�P�N         ��0���P��-���/�������
���� �#�!"#4 B�2B"?!!1xP�O-��� ���������������x^���x@�?bT$c�0!1#AxP0�[�x������x��������h����!�2x�@4�x3BC#2$/xB����x����ݿ�x��������x�!�0A%x0D@311hR!4 �h�/��ݻ�h�ʺ�����h��������h� 2R5Cfx4#334B#!hV2C0 h���ܬ��x��������h��� h!#"3&3UTx$#$3#3#3h3S3!�h�����˺�x��������h����� h$&4EDeEehEV7Tf4F4h4"2���h��̼�˻�h��������h����� !hBDFVFVVhfUETCD3!XD1 �h��������h��������X�� �1C4h3#DCDEEFhEUDSD32"XA" ���h���̺�ɻh�������h!3#$Ch54DEEE4EhDD433"h������h��������h��������h "4D4hFTEdET4Eh34120! h�������h��������X���ݽ���h ""C$hDDDDDDDCXgVT5h��������h˼������X̼��!X"45EFWVgh3D344$3#XcE4" h��������h��������X����  4h""32444Ch4533C##X#��h��������X��������H�����Ceh233C3Ch343$2"1!XA? ����h��������h��������X�� #"BXE%GFEuVeXVUUE4C31X������h��������h��������X ""53EXUUVVGeeeXcUDC22 X������X��ʻ�ʻ�X̽������X !"$3DFXFFFeVeVTXUEC221X �����ۻX��������X������ �X$#%46X5SUTTTDDX3D"2! X������˻X�˫��̬�X�������X33DCEEX5FDDDC43H54A ��X��������X���̼ܼ�X����� �X4%46E5X7D5ECC3AHRQ1 ��X��ݽ����X�ͼ�����H�� #2X2"44$4E4X6$E#D$"#HC#��λX�����̼�Xͽ������H�.1@T65X3335$D$DX2C22A" !H �����X������ͽXξ������X��"#3X$34D3534XB3"#! /H����ͺ̪X��������H�������H!#&U&X3$A443$HSe64#"�X����X��������H������� X !$$X3#$""H4`PC��H��
ܺ˪X��������H���� !X1"!314#X332222"1H  �X��������H�ʽ�ͭ��H���1X2"#$HFTWUF42H4���X��������H��͞���H��� #QHRBbT74FCHsF45BBB2H"���X��������H��������H�� CH4EEF7DdDHTQRR"2H�������H��ܮ����H������,H���4#%X"!2###X$�!H--���޾�H�����ݽ�H������;H2#"BCH44CDD#CHC2! 0  H�������X��������H��� �H QAE44H45C33C!H@$���� H�������H��������H����.H"35CDH3DC35�1#H1�� ��H�������H��������8��+M���%H132AC2H5$@ 8A�.����H��������H�������H�/�H#22A2CD$!���H����H��	���H������H�?04H#33$H!!/=H�������H��߿����H����.H�N0""!2H3$2287"2��H��������8���ګ��8��,���NH!�@"1H$"3^280@_�/��H�����H������8̱���H�21285V1e#3QH�������H��������D������ H��<1�H!�"!2#H1"1�8>>����H�������D����128/0O5�H110!4FDD]��8<\K����H��������D����"DH�O"H!" "!!8C� ���H� ������8������8���-��8N0A1`H1!"!OH��M8��������H������H���08@1 QQ2H 0"?"�?8S .=��8������H�����8����_"HM^0?184!$"H ���8������8���)���H����  8��#�1a08C ��H>= ���H+���4���. "5H��?  8�RD"_P8Q1�?8�+J/.	H�����D�2B8.0��B�08$#RO_Q^83! -0>8/.�á�H�����H�������8��!#!38OU�Q\r8/?��H��,��H�������8 �� .�8�����# 81B?Q1>p=H?���ղ�H�-��D������./8.���n(R�04Q4Q8OB0?]^08!�?�8�У���8�,��
\��D1@Q1BD38�NA  }44�-��8�/ ���8������4�����#8ӵ���"H?�����8�1��8���� ��8߲����4�/B0C8� 0.3�08���O@8�>!��@8ᦰ9��8��Z�4�2U68!�0 OA9����/A�        ���D�_�[ö���� �_���M�O"�3���-�`��.���?�-���R�-��2��^�#��  �A������S�!��#�.�>�Ϻ2�.�>��! ��/�� ��M�r �����o��1˪�$-3�0���V��@�#3������R�E���?���#���0�E������b�/�Ҫ�0�a�ܪ�a�!���=� ?� ��4..��D .���5 2�
��!�C�����@/"�Ҫ$O���!1����O&?����51S����4dݼ�c2λ��3%?��߮�3AD����DT�μ�c3����B%>��ﮚBQD���4t�ݼ        ���L��/�/����1�= #������*��æ-� ,�_���-�����N�[��� ���"S�ͪ� �� A�ı�"��/�� �Zl ��� ���N0�����������@�!�,���.���1⪆�S:�� O���".�՚_ � CD⊾*n�#�Ě��������K��S��!ozc}O2�5��� 4�����N�����=���P1����0��S#b� 10�,���������� ���]�2� @/ �$>0 �C���D����L��/�.��%-����A0����0��D#cҊ 10�,��������         ���R�>���!��S��R��2��A��1��S��Q�.�@�-��C��A��%N��@�?����A��b�Р�#�2��0��6-�B����R�=��E�B���!�.�$�.�" �/��� �O��A��2��$1��W�f��E�A��P�#���!��`�R��`�%0��B��#+�f��4�0����d�# �  �#���Q�� ����C�p��VO��"��"��D��$?�/� ��!��$/ި� 0��e��3�3�"� �D�ѨD��T�0���A��C���F��2���#����_�P���%<�F-��6>�%�E>��""���.�1��!��4�#��P�����e�C����5>��T���"1��$�@��1� ��"�1��#!�����E�,�S�C���5N�a���1��4>���B�1���1��4/��E�>��U/��C�.�2���.��!C�����2����D��E�-�B����1�Ѹ"�1��"���0��e���2�" �?�A�  ��1��2 �1���C��/��D�A����$@���R��3��� �1��4���4��C���$@���.�T�#��U��3Ψ��4�N��c���W�2��$/��T�=� �E,���C�!��2���B��$B���"��C���D�#И$/��V@���D��T���D��#�0��T�!��" ��S��3�����T��6a���D@��3��$ ��&bڬq��#/��d�%� ��3�40���C��v��%0��!���%=�S��2��2��r��2���B�%�D��B��2��1��d��5�.�&P��D���1۱V>���t��"��A��"2숢g.��f-���U-�R��xC�`�x'=�@��Qx��2��! h��#1��S�h��D�%A�h�Q��2�H�51��E.�IB��2�         �^�0�S�Ъ# ���4�2/���2����%B�ͪ32��3�3���#1!����S�ʽ�#2���3�3���3 ����%C�˼         �C ���!��5! ��R���+�C�^������?� �����,���1����e��R��%ɰ��1\�!���]�e����?�# ���1�0�2���2.�"����!��<� ��/"�������%3��� S�����4�"-�4���� B�@�O�1 ���^�D?������5��A��D��1��b��?���,����E���3�^���1 ?���#��3���P�D��3ߨ�N��2��/� <���O��!*�.�# # ̨% !��T����?� ��U��%����"� ��/�T��Ҩ"�2 ���r��$�M���1��0�#� �� /�>�4"ݘ"�%Z����e.���#�S����!� �$A�3����D�2��$Rʿ1����0� ����A���DV��� /��# B��D�����C � �B�����5ݱ?��"
��� U+��.�R��R�P���0� ��P��J�E݈A��&[��S���3��.��c�.��#5��^��_� �G>���?�$�2�� ��$?��/3����D!��0��B��^��& ��O��/� %���=���2��/�2ЈA�Q��/��0� !�3.�� " �݈!�!��!���R���3��A��A�1�A����!���/ ���A� x��G/�괈2���S��/��@�x�FO���#x�C��t�Ecګ��#��"�1���B���Bx��N�2��x.�#O� �t0���T1x��T��x�U��1��Bt-��D�hq�E,�  dA�"3h �#h�1��3�!h��3�� �T$?�"��DD��b���H@�� �48�!�U�"9� 2�"�        z���l�;z�\���z�S�#� �O�@�zM�!W�"-�2��� �A�! ?��?ފ �5.�4��?�� �.��3��������� ۊ/���O���5�E ��%14 �e"c�DT�D�"4?��E /���� �����B�0�������������������.�����!�0�1��E��� � �N��#1�4# "gz$eft3Cֆ���"܊4������/�  �� �����  �� �����F0�"#�P�C��2zUO��f!D��EB""/��d�E�E��$�� ����2���v��U���z���� �2z���b��E���C����� z����@�@�4S��#"$C$B�#2$C0�6�1��4Њ ������������Ί����/��z��%�V�zB �&=��U�"��3�%1��zf?2�#z��-��Cz�  3��z�42��?�4� ��C��3z��C# 6P��%^��B�/�������������@��$1�D#31�B�T �$z#/�%A�7O���������������z�����5�z �G@�uO��#2�!�4"   ��1�T� z""/�2�$z������ ��##D.͊ �0z��B��$Cz $�e�zVd ��R�z� ����z�����z31��"e/�E/D132z#4Ed%dz0�0�D1zۼ�-��۾���������z�ڪ���/�����4/�zGP�R��32�#�1%T �"z42 V0�z������z�������3��z������4/j���5Q��C� z�����z���ʽz4?�3wzS"DUFVTE�23 31� 1 �3z������z��ʫ���z�ˬ̫� �z�/��D!!jf2Vs��"D�2� #C2!zCB W11z������������ ��z��Aٟz/��4��zEB�!!�z������zۼ���˫�z0��2��4�"!#24B�"132 z5UR��5C!z"B���z�����z��ʜ���z2��#?�zE1�B�# z��fS�Tz�%f1$VzT3#Tjc����z��1��z��3��4/�z�����z@��A� z"E �"2 z ����̊������z����Uz?�EB%T3z5U �%T0z6T ��Tz�3 �� ��z���˫�۽z޹��ܫ��z!ʿ"�3jSB2CUuz�ET$T��!!$2z3C"C3"3jb%B�ۚ�  �� �z��!��z������"z ��#��z3"3!j"�4��z��.���z��50��#"z"2$DB#EzfR"4Cz$eA�C �z"1���z����ܫ�݊��������z2�����z!�!$Rz�E1��EBz�"!DEzU2#31C3jDgB"F>��zܽB��j����z��! ���j.��4A���j �Ec�Ez! �" �z�����z��!�� z"#3""5ze333EAz5C2!"!jGP�4��z����ܻ���������z��������z!"�E2�j�e�fBz��E2z"TS!"3#z4A$C/��z!/��!!��j����z�����j-��d/��j��Wr�tj2$�f?�z������z�����z4#"6zTC2D5AzD3B"!jG`�4 ��z��������������z��� ����z"�DB�k�V �$fQ        ���/ � Ϣ@�����#��=��?�<���2�3�����#���!�@�E�n�1 ��-�#3̢���3d#ϲ���!���C2����"?B��Ṟ2ݪQ��S������������aN�B/�!���3���U۲lϺ �=߶�?��O�0�2��B�� �.�O�����$o�����P,2������� �=���=�$"B���.@^���0�  ������2������.�C��.��4���� ���C2�V��M���� ��У&Q�����3        z��C!��j��<���z / �!�!�2!j;��� ��j�� ��d!� 
�RjU̻�P�#j�������jCDC���# j�E���z� ����d� �� ��C�� � j�  ����z��'5B�"� �@�j�_/� <�� ���B1�  ��0�#=� �j�����͊�42�!��2   j+�P �ݚ � �2!�  �!� z"[�� �  �  ܚ! � ��#�D!��j�_�!���  ��Q�    ��0�O��!� �    ���4A �/�3���s��j*�1��� ��!"��  �A z��!�/�  �zGTA�� ��?�D�z�/  �5���@ !��� �$ zB���  �#�22 ��"���A � �    ��@  ���  �Ez�/  !�  �2  �B� C��D�    �Ӛ`���� �0�C!�j_���D4;��2 � ��   ��B   �   ��?��1�� � �  z 2$��B ������몬� DE�  ��!����C � �  �1  �""3B5~��A ��  �,���#!� � ���!2"�� �#   �    �������$�  ��Bz��� 0� �  ��D ����0���  �@�!���#C�   ��� zo�0�� ���EA���C � �� ��Q�����"4A�  ��A z4��$:��$ ����E0 �&�� �����1 ������#U �  �S ��! ��R������ � �o���33� !�  ������%C"�   �  ����"�Qz��/�۫�� �����""4C"� � ������D#2� ��! �0��@ ��������    ��S.�   ��6 �������B4� �2�  ��?�;�a ��!�����   �0�s���U �,� ������D4OѺ��    ��d��A��z/������  �C ���  ��D���"�������5c���1 �  ��1/�-�za������""4�zRZ���f�1���̚�� $/M��B �    ��"��!z��������0 ���" ��<� ����� �""4
���4VweD1�-�� �������7�#B� �2��A�"�����ݶ ��#-��TS!�Ί! �,� ��� ��@��3  �N��3�� ����� �0�Ee!���!�����  ��0'�#�!  ���$�/�+z�A���!޶   1� ���  �1��#�� ��6�R��#DDC�N! 1�N�zQ�����   �3  ��.?��1� �-� ��ަ�� �L��P �� ��#�!� z�� �.ĺ  �4  z�q�14�^z�J�1���      ҦDD!��z_�"z���@�L� �  z=�!A�zN�1!���     �@�C+��.��za���j��+&%�\���   ���� z�""���R�    �A �q��?�2v�@�����j�M�c�[�S��$ �� �ڽ� ��z�3��E�   �A����$�j~���$R��     �" ���zW�/E�=��zC.��1#�  �1 �z&���~��]z��B���   �&�c4/����z�V�P��#z ��@���B ��!��0�_z�A ���  �4�3P����z`�!Q�� �  � �C���A� ��� � �z!�B���  �4 za_��2��@� �  "��@    ���/!�%z�B�!!� �C �Q� #��E  �    �Úb����  �"�z"�2��R � �-�� ��S �  ��?��1� � � � z�C5��B� � � ������#34� ��� ����C��   �b �#3CF~��B  ��� �  +����##� � ���!2"���6 �    ��������$�  ��Az�4�!0� � ����D ����0 �����0������#C�     ��C3"!3#��  ��DB�         �b��$P���"��S��#�>�# ��"�@��#2��5�O��1����E0��5-���f��@���d���D�.��%P� ���D/��     �#���$��2����GP��d���V��5P���2�� ����e �S��%C��51���#?�!��3!�#����&�P���E/�ި�V ��U-���2#��#�#0��C/̸� �/��S���3�Ш4U��%R���D��#�B��$C�θ�/��C!����3!���E@��4 ݨ� %P��4�?��C�߸"��3!���DB��#�C���#1���$B���$1�ʽ�F@����1��1��4"��""�-��#C�R���!����#2���T�E�јE4��"D/���#0����B���"�����4��4!��"�C ��40ݘ�"!��u����C���5��4 ��"!�0��31�Θ!��g,���D����#.͘Q�C!��� #B��"��V.߈�W.���"� �/��b�33���3���3�P� ��&O��0� � ��1�/��"4.͈�WP����# ��R����Q��� � �!��2 �0��"$ �ވ�4S���5�2��C��D���C���3��3 ���#1����$D?���U��5� #��� $@����U
�E ��"1����$0���EM��>��#����3B�5,�5! �ψ#%D����U�"��5^��0� #����C��=�40��45���D2����5O��_���FO���3��&+��$0���4��33����#1�P����5C��ވ2"���FS/ۼ"D� ���#2���A�A܈��4C���x%5R����6�D ���#2!x��DD/܈�� 4/��x�6eBʾx"E1���24xA���!3h̜�%T/��x��V@���h�VV/˫�3i%a��!�         �� !�"Ѐ�@�G+�P̐�/�M����O�&�@����0����-�����?�2��   ���g���D��O���A0��-�B�� �p��g>������%0�!ބ#�@�" /�/�4��M�A�$����B��4B���O�1.�^�2��@�P��@��Q�1�Dݰ$��-�@�2��"����O�Д.�O�0�/������"�N�Π �O�c�TݐV
����� ����"��?�U����>�}��,�1���!�� �NB��"�!�1��?��0���!�C���� C�Q��ڤA�@�=���@�!� �/���,$��#��R�� �1� �<���?��L����T�]/����Q�?�"�/�?�.��3�O����� �"���2�"�����Q5L�Τ-�� �_�6������@��G��ѻ,W��V�>.���@��-� B����^��C�^����� �o.���2����/�1�a�!���Ҥ, ��>�� �,�ң�\��>�����0�Dװ���� !�� O�� ����!�Ұ.,���1������� ]��;#��- �����-!���2��N.��KP��n>.�����_ ������/1����� "-����4���.�������/� >O> � �F����N��>!����//��� ,��/�0�..����q�` ���6�����ѐj& <O������1����  ��+@����_��B�����.��0�߰�!�R�-0��� ����[���.����] ��]���!��>��\�3�=[��
���=���P���OҠ�ZC��-���?� ��!�/�����%��c����N�-4�.�.���
����1�#!������"��������"���� ���=ҰD�c�1���?���1,�!��U��b��%� � T��F�41�Q�"ߘl�NB���x�1��t�Tb���" h��-�Y����         �A��@�1����0����_�3���?�����#��"�^�B� �#�!�6��"��z�f��O�� ��@��#�0�C���/�#L�R�#2�����RA��;"S��Ԥ9"���ߤ� �T1��̼��!���  @��!!����t��Τ�����S1 � � �� ��   A¤$CZ�����  �AѴ$� �������' $2�C!����x^����@����:�]%�/�^$��3.�ETܤ���$@�������.� �Q� �2�!��� ��DD1S�����T�!"��ܺ���N5dB�ۣ�Z������"$���������"""��}�U2٘> !O:���C��1� ��>�<!����@�!>��2���p�6� �1��3��  ����ED2àd��D1#ET�����"! �*"����Ш*6�� � J ����4!����"���A""���3��
��E3����      �������DR$�/��/ ������DD1��<�1 �+���;��C����l��A��������34Ux��� e"0� �@��� ������?�?x������Sxw���� x�"����Rx 4�C1 ��� ���� �C�� ����/���  �����PS ���� TfR" � ��?�������� .�A�"�@�� ��  �KC���.Ѹ��� Τ>D�����1� "�����!��1� ��+ >� ��2<�&�4���o�1� ���3����j��  ���@��_�##�˼��"$4� �
m���D�P�<�/�!��O  ��=0�h"nTR�� ���m� �C� � �@��E��A�������S �=,C[�  ��?������ �0x1��0R3�  � ��xL�3!V�ޔ�����+���   �������3�"��C�?�Tߔ$��>�O�!������>��%5-�"3��N2;���/ � ��0��3t>�/��64�p� +��tb��� #E�  ��O�!� ��4,.=���"�1 �"/���t2�,� d;���a"1t . �h�    TQP� ���(A� �8 �����ۿ� 4�4  "#����          �  ��$] =��p�B��Ԓ��������O/ 1�Ӗ��NԖ�� 0����� ܿ���0:�RӖ&���1o0����2/������A �4���@!>��"�!�?�R��%���`��P��&-���A�B� �5�.$���`�>�#�U����O�_�/�T��T���~ҶB���0��M�n�N�e��#���N�B���0��/�?�/�3��#���?�C���1         ��l�;�˴��2.> �����ߤL!#S���� >�Y�Q1��������0!/1Ӵ�O�����������!��/����!0S�Q�?�1�0��AC/�<"S �� �0�?��%��dN�0Q� /�-?,�����Ӱ���T#�$�ݾ �?�,`�1�������.���o�=�����0��Q,$?��:@�"���2!3 �B  �2/���3� 2�����3�o�,�����/�0��Z!����ԑ%�O�_P�L&��U$AE�=�����E�$�#�A���@�,����.�<��-��C��5�0�!�B/3/C�C�n%#��/�_��-!�����O�/�����A���!"���N��B\�O *���[�/�_�Z��
�#�0���\-�/�,�Q���]���������2 ���? .����0ް/����
ð��T?b�a��.�/�,����Ԯմ����m������@�"�$D��/A�B= ����F����
�?>�_�L+! ?���������P@B<�Q >�?��2�^�"��ĥ���O�?S5C$���/�,L�=20�"�a /��Ӱ����0��.�M��������N�>�-�A�0@�������д�=MM�M��=N@� !� ��C�5!�O�N�Q���C@��!�/��a�0�?�����������>�<�=��.DD��;�.���M��0��B6O!�1߰B�@��.���A�/� �\��=�35�#+��2�C"�4��D��?��A���mN�@�1������ ��3� ����Q�=а@$B1�� �C!�#�� ���,1��-1��K��������VD_������/�M ]��Y�J!.�?�?�@�>�߰��/�[�<-l0m���Q�&�o��"�!3  ��/�_=��0�����������?�#"v35���.��,���"��Z�[��>0$����#���N�<��--����3�����������/O� >-R�!� �� ����-��Ġ��R.<�� �,���٠�C�@>���������@�.����!��<��& E��O�0.��-��"Π_�>�����3�A��� �!�%4�C�P��>�- �������- ����������� �" ��?�
<����� /ސ$� ��2ഠ��2/�/�A�EF�����.!-^��������RF�A�>��.�J�M=� $�����/����!������#�� @�l�9P�a�#�Ns�N�T�<���ɠ�"���`�R@�1��>�%�?�5� �1��L!�=��!�$�"�����۔/�L=��`����"��3�1a$-�#<^�����T�ίN��߀/2;1C�d�BU��������1��1�]�/���.��B�!�A����1�/��o�-K2�W�$�U� Ӕ+ A�S��"�!�/�>�33��N�o�=K��!�0�M� -������p��
 ��A� � �-���� �!��2�!�<����$��O���+>3�1 ��������QB�"P 1�� �>��O��p �;����p�������p�����p����pѐ�1�/�p>CL4?%$p ��.�?pA:���p%��.�Qt+L��4�p����"�p?�.�
>4p�%$�4�.p�  +�- �p�������` ?#!O�`�.� $�`4��A��p1��p� ��.p!B �"�`��@� `�%� �2�d�1=�Tm���#�ud����`� ���P�1:_bP�t1r�d+P�0�����P0�>�_�P����P,>> �T������1P� .��?@�@�E�@Tq�.N�@.���"4�,�\aJ�-4 /"�Q�0������0���  4������$+R.0�?$�� ���$.  ���� $ 1B �?,��� "�� �0�  �0                                 �1  �z$������z��B �C�   �{4.������         ��N�:J ���� "��2�P�0䖰vRdPp#�"�,0?����� � ���-5����? �_� �+,_�� P��� �<ݯ����������@/R�7ִ� ���..�+�V��墴/��M��*�������O�E�+�o �__� ��MP!��n
C��2ߤ�Ҽ ����Ӷ�? �2��<.�jn���N�;��- ��.��?���������ձ�ѲZ�/-��.�/D/�A��n��4�QM͠����ޤ�/�� ���.�.��.���� ��  �Ф��-��"������ ��&¤��!��"�AA����O �?�4��"���/>���������?�M�;B�23D$32�=nZZ$��E�@Eϐ3/"�����*E
��0R�TBM�"BO�=��@\��T~���2����ۿ�]N��1� �A������!�͐M-n����]D%��fE������;P�0@� [��\�L���!.�,��2`��R���N�N�=���42�_U""@a����0��-�>���A��"�N=���C /�A �0=ߔ�].� 1ѐ�1�/DB�  -�0�-��--O�O�.�&�-�DM������23�/ �� �-���� 0<O>�0M�� � �����]��,�P�l��]m�� �/"��c`B�����������$�D�0τ���n��$�23?!߄��k�6���C$dF4WT�%�����Ѐ�/�3��]���t�1">�>�EcR�=O������� �������
�#�EU�D�S�/�!?��2���B ھ��# ��41���� ���"���t�q��@It������@p��
��$Tt���`�-�1/"�tѧO��K#����-/tL!��.��p ��dt�l�N��pS�Qڽ���d�o�[ @p ���)�Bt/����"t� <�.+�t��C�=�p#�C2�tB �!���=`������`"�U��TGt"�, �t����p� � �`�S�#$PTd�4���[�d��Ak�d �/2��d���1�0d �."��0�d� ��,�d��=��L` ��P��D"-+-`$�-��PA,�K,�T�I6��@�QP���P � 0T%1Ed/���T�PO��2�P3� 4?2T�N�B� \�P������P�?�P #13O�P/������P��� ����D���o��PVT"�D4@�P�P�D���q+�4���n*/D���"���@����,��D ����N�/4N�,<�D�+1�.�4> >�B�-�0 5��� Q��!4@����4 ?��$`�<�A�$��- ��- �/�S�  ! 3 _��n���k�@/��� . ��
� �  ! @ �      ��         �                                          ������   z��?��1�  @�!� z�f���{��?� �1        jDd"�z �����z������z��$C�ze?�%fT��"4B��!j�����z����TBz�� �!z���#E?��D2��z2���!z�ɮz˯��$R����C�ފEA���zB"���ez1����Gdz��1�C0����%T��4T0��zB�ۮ � ����z�����e>�ۼ�EA���E3�� �!z� ���������""� ��5c���5T �$�E32� z2�̪��!�˼� �� ��ER���UB�3zvS3!�  ������ܻ������!���5f/ފ�$T #3zfED!  ��������� ��� ���Ee ދ�5C!C         ��R/��O��^�Q���O��߀�c���Q?�ڼR��"p���@]�ހP>����?/� ���! ��/�B�є��?A철�#1��1�A1���"�<�M��ˤ���/ =�� �B!-�3� ��?1 ���"!�D��4.��?��+���������O�"!�k���1�2��!��"�������Ѱ�4�����!��������{� ,?Y\�a0��" ���   .N�>��N��@1� 0 �nB��p_��?-��   �����;]>. �^��=�Am�,?����NO� `��0����    ��������p������Q?�?p-�"��ZN`�c��2� �N���@Z*O@���!��2��1/� !>p1���"�  �"�5�L��A ���/��2��"�@��E��1��?00��a����M���0��@^�!�L^.;AeC� ��!�D�# �L � �K��� ��� �C/���3��"_��#?��4͐�D�_��, %���&���!ݲ�"������^ #��  �9���> ��.��Q�B�����"?���A��U/ʔ�S0�D�� �4���Q��!�����B����^���"�@�d�.��O��B����>�.3�_������P���� �<��R��C�����D@��#��.!���  ���!��$.�c��*�2���P�4����/������0����C>��0.�O��N�? ��6�/� �� �P��2���b��C����^�,�$ �!!����K��Q����~��ԭ/��" �� � �$,����2����2��.�����P�;��UK���      ���E�B��.д� �e�_�4� ��R��/�� P�$N���]��� �0�#�5`��"�#/��_��d�>��� �C�!�F�0�B�,�?� �d���E ��"���C��A��c�� ���Q��3� �!�#�#N��  �M����@��2��D�'=���E��S�23�$�=��C��?t� q��1��,� �3���D� �p�/�!�p,��2���tP��A��5t��] �@p�� ��2p�0�����  �#�2��P� � t� �@��$t<�1 �0p� #�`#����5�/�           ����2Q��̿PB �O�� �2�A	��O�1����22�� >��1���4"41��2 !��������aS>��a2�-ݭ��R?�޿��R2!@��ψ�5��?�/%C�����T/�� MxY�����m>"A�..�����4�E�Ϊ�Pd�A�������&����">՘b�����5�?����a� ���3/�5^�-� ��%# �����g/���� �v!阺�LUQ�����"Q>ʘ  �!�' ����1>�-������.!a�$� ����S���0�6/����7;�Q��_��AΘ�#��� ��R��3� ��!� ��1���a/�Q�����D���  ��� 3�θ��2�?���� ��� "����._@�]���3 ��<��_�"2����%=�"��/��3����ScE�̸���<���D�3�� ��C!�\����?ҘN�.�a� �0�1�5.���# �!�/�"3����^ L��	�?����?�/�2_�O����������3?��C���#���B2����o, �����A�! ��Q�!�
n��ߟU��T#N���T��� U�Ψ�3�->���o��� !�R ��#!��13�о"���R��"�?�A ɨ�c"��S�!?��1�!�.� U-���!� �N��N�������D�����#/��0��!�/ݭ$bܨ�S���&� ��`*����3���#�� 1.��C??��#!���2 /��AQ��r����S/�/�C!��f����Q���5��  ��2
�T�^y�F����11         �������̸  ��@�  $���� � #=�� ��� ��DC �����@��M�@���=��"���332���:���5B����o2���&��.�[���b����!Z����!/���O��/��A�-���[���/�0������ *���/3���%0��!�N�?�ޱ�0C�!��!$>�b4_���$� ��4��1�0��� ��.�M.��N����P�¸O�/������N��,0Oϸ?��$���?��"U>��_�C;1챤#�1%�.Ϩ���@��<��A�%�-Ө �Z�N��$ ʹ!>���0#�`�� ���_�&�^�����5��� ��B5�/���1� �����D�2��a��޴_��3����-�$N�1��1��!�5 ����CL���aޠ"�?���!�.�^�+��F2����0�1���-�01���  �.��!�@!��!�B#�!�  �N��#Q����.����3 ,�/��B�?��!6E
��/2C� ��� 20��=�� tΔ�˧OW����$RQ���?!�N���e#�3����^����3�� �#B��� �E�l��0�@��-�A�o��� ��������K� ��?��03>��2��"ܔự CN͐����ϐTO��S ���A�6�2�@�m��C-���"��"#��Ĩ� �.�O�/�-�+%��2�0�Bϔ�N%�U٤�/�-Р�! �$�����S2!�� #?�ܘp`���"��.���4!O,���?k�^?��� 1�ܘs�R�0�B���<����"����"-� ��+D��� q��.�23����/�0//���2���� 3����#����1���R��# �"�����=��-�P��R��f����QИ-�! �1����`�#GL�����N� �1�"�?�2ӈ��@� T�����N���>���-�O���B1���M�\N�<܈B/����� 4�=��O����=�4@@��fO�� ��1���1&�!����O�$����E��5/�"	�-�QK՘�O��2��R��"�+���1�2�����!b�+��M�d�U���>�� ��$�#�1�/� �/���D2����1 "��.�2��@��C���B"��%-�?��W�1�!�m����F�N�Q�$��&����!���R΄,��S3��2��n�s���?��/�" �?���M�#
π�� ��!  x.�\���tDC���b�1���b�P�����S܈ ��d!���O�����- 1�x�^�@�N�>x�?O�+ ���$A$=�ވ�c��)� /�-��A"߈^��,"t�"U! ��xq� �}�x��/�R�$x=%� �!x�>�4��"����3@��� �e��!��D� � �xP�^�-��xBC��Mx-����xc>�\�/�x@���O�� ���x -"���n3x��+�A�x�$�3����#"E,��@È.2� �@���0�31��x�R�!��;��!�%O�/̈1�D�=����1  �x�R�=�t� #4<��x ��/�B�t`�"��-�x_���0�%x�>�C�.h� 3�b�h��1?�h��!��h�P"�� d�"��$h2�"��T_�#-���5X�,�R�CH-��<�UH��#�2�8P���4(� ��B�S)�!��         ���?J��Ђ..�"�o�M��j��q�n�-!�� �\�B������r�!� ���3�ݦ��C$���O=�=?�ѿ��2�����%N2���/1��>��D5P��,'!R/����pAG;�����=c��c��𱼆�U <���!�$N����Q�����#D6����/A �ޝ�R :�����"����N���#�����#^ Q����J�l��1� 4B���! �� � �?����R����C1�ۆB�N��d���$/��1U�3�/���$..� �v@"@���r�� 6bB��!�>�=�_������/!!��.�v�W+��#�v��/R ξer!�C! ��r�D��"!r����TN���7b����C���3�=����/��A�rb���"%r���2D ���M�v2<@�����1 ���`��1��K��?�B �L� 3��3��T=��@�"o�� ���O!� .���4�� ��#�3 ��E_����b��E۲2��&=��5��/���b���< � !!����6���$.� �  �@ ��p &���2��"����5���� /" ��� ���N�!������� � �ߒE� A��1� �����PM����./��� ;�� ��K�\�2!�!O���.1���ϖ3�#= �r��5A	���D�� ��b��?�0�2�"�b�1� �!�,��A�M���#��0�Y�1�O� ��lѠ?�?����T���Q���D�^���3�3�� �*�!����$2 ��1r���3#<�$r ?�SA �rT��$,�M�rB�"N�F܂#�2�Q�B�r��/�'1��!!��3����?K����������������               /z �L$��/�� ��2�U��Pa�� ��1��2��a�ӪC��S�R���S��"��c�� !�Q߬"�B���!Aޭ"��S��#�1�!S����# ��B��3� �!1���#!���!@��3�0��"%R����# !� �GAʱT �B���7B���T 2����6A��D�2���FQ���3 2��ܚ�T2 ��B�"���V0���C�ݚD!/��2�#����D ���"""��ܚ�F/ ��2�3����4 ��2 1����#� � �1����$��"0��܊�F��5�2����4��32�D�$!�C���$� �#"1 �ڊ��!  �  �� ��A�ي��&�1!������$ 1ˊ��$�  ����!3�z���/7"��� z#=D"�z��63� /��"� # �z���5D��  ������" �z�D���%C��� ��" �z�!��/�5Bz���"��z#1#�z�@��$Rz"��A�ߊ!! �z�O��%Rz#��0��{�R"��        :�4#�� J��!1�ZO� !�J�&���Z���T"��Z�1 !Z #1#<j���4e!�j��2" ��Z3�?�"z����%d�j��D!!�j4�%A��� 5R��j��BV0�z���ފ���W@��j�b$A� j3U!뻊 �%A��v?��#4D2j"�܊��� a��� j1$B"!��  �r����  Z���������A����!�j� EVD/��   �B�ݽ�  j������ � ���$�B��� z@� 3""� �����C��� ��� ��� ����듪T�� zA� �3U����۠�F.�� z�����"3���� "���A��  �5B!��$z2ܽ��۪�4/�� jVk�����B��2��GO��vFUT!��z4 �� �ʪ�4/�� z5-�����!���C/˚�F?��!jQ$ ��$Vz4 ����ʪ�4/�� zU-���� ����3/��GN��v�eC"��%z3!�� �ʪ�4/��j������4���� ���V>��jVA� �fz40����ɪ�4/�� j�& ���Dz"˩�۽��WN���!v�4D2��6z30����ʪ�3/��z����"�������4/�� zQR�  4zD �� �ʪ�$ ��zr� ���"�������4/��z�  4zD!�� �ʪ�4��zA`��$������ͪ�5 ��� v�!����&z31���ڪ�3/��z%�� �"�����˪�#0��� j�R"�%gzC0����ʪ�4/�� zB� �"�����˪�#0��� j�b gzD ����ʪ�4/��jr ��E�����˪�$0��  vb��̻�zD ���˫�4��         z�_��4�zs:�3B;�4z���6���bz�.�C ��zc.�f��az-��/���� P��M�0� �jQ/^�U��~z��$��b�z�V�#ߊ�1��1���!�#�1��S�z�0��#���2��1��1���@���A�D�/͆�n�S˾$D�=�C�/�A�T��1��C-�E/�����51����e��1ۚ0���-�T����B�ފ5a��B;��2�<�S��C���2���C��d���1��1����s�z2�5�6�NzWL���Q֊,� � 2��M��N��T���t�Ίn�/��  ��1�����Q���5=��2�/�j��a� �2��!�Q���"���Q� ��!��2ߖ��/�2��B�#?��3/�D���
�4
3����&�e�"�� ��%�$��T��M�!����%�?����B�� ��!�5��0��T���  ����c��%:��� 6u�ۊ�!�6���M��S��q��#���z#�O%�!���" ��D1 �/��A�����2�2���$@��3 ��?���Q�1����f�� ��! ��1�2��#>��C����4.���#�,���D_�� ����A̚1��13��@�� �Oܭ#?����e���b��1����1�0��E�	�"���G���5�!��Ҋk� B��+��@� ��C�� ���3!��3��b߼""��.�  ���A����B����r��Q����6>��.��L��5�@��F`ЊA��/O���A�� ��-� �#"݊�6>�G ��"3���0� �"���4@���Q�$T�����!��d/�E���S���P���0��D/݆�m�gA۽��$���Q��3��c � ��6@�����?��S��2��?�z���l��� 2�1� ��gߚ� #��4�� �$���� �����$ �ޚ2!��d���#��"���#2��"�-���ݚ�!��C���D����C���@���B��P��%P�#!������p��5�/���b���$ �-����$ ��B��3 ��?�����L�!���P��� �U��$��!����C�1���!�����1�1͖�d! ۼ�����3�!"0ݖ1���ݚ�"�1���B�Q�0�!�7<��?�.�A�����O�c���3?��2���$ �>Ϛ�$� ����Q���c���@���D.��"��4��4.����B�� � �4�1����S����1��W+��O��%-��0��s��# ��}��@�3��ߚ ��$"��1 ".��$����B��"�#��6-�B�����3�!��?���B�ߊ�p�"�ҊE��6��%�A���c���2rQ�F�^ܭ6A�F.���.�^�A �@U.��s���5�>݊2D@����"3��ϊU���=�  � ���S�˽�d�!��"�2/���V0컽�\�_���!�/����A��A�К?��! 1���5?���3>��-ފ�!/���$?�/�����N�?�� E=������ߊ���0 ����U.��� ��ߚ #3���U� "����>�"���Q�T�� ��/���4�Ϛ Q� "������-�0��!0 ��B�������"C@Κ�D/��A�� ����,�!�� � !�@�.ϊ&O��.���3Ί�"��� ������2���$/��/��f�-��FC�;�"����0��" �.��D����E�$���O�����2!�@����2�њ!3��B��N��R�����2 ����b ���F�=��2�B���!�3��C�?�$��2����/�� �̚�C��� ���#��5� Ú�@��$�1 �!��A��"��1��2 ���s��$����31���D  ���� �!"���1��B�4� ��B��!��C����D�?�"����$����1���2"�?���B ��A�B��1����"� ��#1�^��Ba��/��A �� D���d���N���Q� ��G��V� �5�C���5���?��!� ���E��@ �E#������"�"��T���0�� � ��D����RA�� ��"욡S$>�"��S�������~��?�T?�4�5M���Q$�/��1�/��R��0�0���������.�B ��eW�,�#�$�20���G@���]�o���
����B���S"����a��!��S��W>����>�C̊2��?�/Κ#!��r � ��#0� �2��O��f�*�3��?����_�>�Oњ��2 ��A��3/ޚ"���-��3�� ��]�������$Κ2"��u��B� #���3R�#-���0�������$���B���D����%2���O�2��$?��U��6_� ����@���0 ���b����3/ ��� ���1��C ��O���0���L�!��  �Q����e�-��=��0�?�.��������!�-���u2�����%��4�!�"1ܚC�� ���"��2���C/ ��R�?�1�&=�"�?Қ.�@�����0�c��D/��B ���5?�>Ϛ�$�  ���Q���S,���Q���E��3��3.����C��� �D�@����D��� �0��W:��@��$-��O��c��" ��n��O��4���� $"��A�!=��4�� /���1��"���E��B���# ��"v�!��?�!���2�,���`��Қ"�����C���c���1sP�
E� ��!���.�O�1�@U.��s��4��>͊2DO����"3�� ϊd��>�!� � ��c�ۼ�d�!"��3 ! ���gs���$�<�P����"� ���������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                � �0�@�P�� �  `ЏХ���      %�gыѢѦ�      ���*�O�uқ���  ���#�T�nӛ�    �������3�^�    ��������  ��Z((��<��`}��P���F��T�� ��<�Ƞ��`}���T����d��
`�����}�K�}�K�}�K�}�K�}�K�}�K�{�I�G�E���d�  �`��ȴ�}�K�}�K�}�K�}�K�}�K�}�K�{�I�G�E���<��`���x��}�K�}�K�}�K�}�K�}�K�}�K�{�I�G�E��P�F`}��T���P�<`��T�� �P`}�T���P`�T��������<��x�}�K�}�K�}�K�}�K�}�K�}�K�}�K�I�w��<��x}�K�}�K�}�K�}�K�}�K�}�K�}�K�I�G���P`}������� �d���`}���M�}�M�}�M�}�M����d���}�K�}�K�}�K�}�K�`}��0�����d���}�K�}�K�}�K�}�K�`}��0�������`����}�{��y�}�{��y�}�{��y����`�����}�{��y�}�{��y�}�{��y��<��x�}�K�}�K�}�K�}�K�`}��0���*���`}���� �w���y�����{���}�����w���y�����{���}������$�ɤ��y����ɫ����w����w���y����ɨ����w��ɡ��y����ɨ����w�������w���y����ɤ����w��ɝ��y����ɤ����w���<�ɤ��y����ɫ����w��`}���� �w���y�����{���}�����w���y�����{��������$�ɨ���������������w���y����ɦ����w��ɣ��y��������{�����w���y����ɣ����w��ɟ��y����������w���<�ɨ�������������� �d���}�K�}�K�}�K�}�K�}�K�}�K�}�K�I�G� �d�ȴ}�K�}�K�}�K�}�K�}�K�}�K�}�K�I�G� }�M�}�M�}�M�}�M� �w���y����ɫ����w�� �w���y����ɫ����w�� ^�n�� T�  ~չ�������*�  J�X�w�{�֜���  ����x�`��%��  ��(���������`xo�]��o�]��o�]� ������������������
�$���ȓ��$���ȓ�������o�]��o�]��o�]����o�]��o�]��o�]����
��$���ȓ��$���ȓ������� ��.��`x�o��`�o�]��o�]��o�]� ��������
�$���Ȗ��$���Ȗ���o�]��o�]��o�]��o�o�]��o�]��o�]����
��$���Ȗ��$���Ȗ���.� o�]��o�]��o�]� _�M��_�M��_�M� _�M��_�M��_�M� �;��;���7�?�7��;��;��;���7��7��;� o�]��o�]��o�]� _�M��_�M��_�M� _�M��_�M��_�M� -��-�m�g�o�-��-�m�o�-��-�m� ����/�����/�����/�����/� �z�y�?��x�v�x�
�v�w�y��0�x��w�x�y��w�t�x��y��x�w�#x� �I�Y�I�y���Y���i�y� y���0Y�y���$Y�+�� `�� ������������ ������� �������� � ���� ��  0�=�\�gف�  ��  ��������     �  �#�/�9�W�  a�  oڇڑڛڦ�  ��  ��������
�  �  *�              .�J�Xۃۤ�  �ۿ��������^�� �}�0�$��$���0�.���$��� }����������]�}��]�}����0����`���]����]�0��m����`�������	��0��0}���ɲ��D��< �	��0��}���ȷ��ȷ����`��
��0�������	��0��0]�����.���	��0�0]�����0�����$����}��� �%��0������������	�����]�}��]�}�������	����`��8���}��
��$}���$���$���$��� 0]����������������`����0]�$�0M���������}���ɴ��ɷ��ɻ.��$}���$���$���^� 0]������������������0]�$��0�$��0�$��}����0M������`��}���ɼ��ɾ$�
������� �����$����
0����}��� �%�`��0��� }����������������������������� ����	�����]�}��]�}��`������	����`���8�`���}��
�`������
�}��������������_� �$]���}�$]��m� ��� �0}��]�}�$�� M��0���0���0�  }������ }�0�$��$���0�� �	���]����]�0��m�0�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 �T�z(�(    L&'                                                                                                                  �    �                ��G�������� �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � � � � � � � �           � � � � � � � �      A � �      � � � � � � C       � @      � � � | � � � �  c !   @      � � 1 # � G  |� � �            � � � � � �  <                � � � �  ? � � � �������������    ������������               �                        ?              � ��3�������      ??������   � � ���������        ��������                                                                                                              � � � � � � � �                  8 p �             p g � p  �      � p        8      z � �  8                                               � �   x a �       0 x � � �  � �  0 x � � �    X �      �    [ �  �������������?����������������� ��x�����������  xx������������0� �????��������	����������������8�8�8�p�������������������     � � ������          ������  ?00�z�f�    ???? � �������������    ������������ � ���'�8�g�/       ? ? � � � � ��� � � � �     � � � �       �����             � �����~�~        � � � ����6���6� 9 0   ��   �<�~�>�� ���  � �  ?    ��?��A�c�?`8�������������������������������������������                ��?��������    ??�������� ��6�>���������????��������q���� 7`a����������������~�����C�G��������������������W���� � � �����������������������������������������������ρ������������������������o������� � � � � � � � ��������� �`�`�� � � � � � � � �    ?.�.��         ?  6�1�g�'�?����  � �  ? ? � � ���0�� � � �    � � � � � � � � � �             ?  � � � � � �>          �����������������#i`���������������������                 ��������~��� ���������  �� ������������������������A�$�|'���������������������� �!�c ���    ����������������'�#�m���   ������������������?�h8�0�`�`   �����������������@�@|�\������������������1s{ x 0        � � � � � � � ��8�8�8� p p `    � � � � � � � ��@'� �v v r `    � � � � � � � �� @�G g � `      � � � � � � � ���?pq� � � � � ���>>  	y � � � � � ���   	����.;�l�~�w��H�<   �      � � ��;�3�wX��|�~p��   8 X     p �                               �<�����    ??����x�8�<�<�8�x������������������ � �           ����������������          ?                        � � � �                ���<�x������������������������<�|�������������������                 � � � � � � � �                 � � � � � � � � 		  � ���� � � � xp��������x� � � ���        ���� � � � ��� �        &2 p � � � � �          � � � � � � � �? ? ?     =  � � � � � � � � ?���>�>�  ????������(�������������������� � �Ќ � � � � ����������������                ����������������?�?�0�p�`�����??????���������������8�8������������������</?�!�7������������������<�|�x�����������������������;�l�~�w��H�<   �      � � �          � � � � � � � �        ?                 �`�0�0          ``0088 ��������������  ����������1�(� �$�,�>�B���????????��  8 >731         0� ~ < | � � � �00      w�|``000� �  ����������88  �F� �  � �??          ��������������pp!  � �N�.�<�L���İ��88    � � �      ?c��A� �     99qqAA��������   �������� ��� �`�`_���� � � � � � � � �-�!�p�0�O��3��  ? ?  ?  � � �  < ~ ~ �8�8�8�  88888888 s1�{�{����w�              ��`� � �` � σL                 ?   � ��?<<        �� ~ � � � � � � �8800      <<<<    � �gc1         88��/�g�s�/���     ``p      �p�p������t�p�     ���     � � � �� ��         � �  ? ��	��        ��0���o�?�Oy�{� � � � � � �    ��0 � � �@���?         � x <  �                       � � ���0�3�         ? ?���&�<�$��8�    � � � � ���?pq� � � � � ���>>  	y                                               � � � � � � � �           � � � � � � � �      A � �      � � � � � � C       � @      � � � | � � � �  c !   @      � � 1 # � G  |� � �            � � � � � �  <                � � � �  ? � � � �������������    ������������               �                        ?              � ��3�������      ??������   � � ���������        ��������                                                                                                              � � � � � � � �                  8 p �             p g � p  �      � p        8      z � �  8                                               � �   x a �       0 x � � �  � �  0 x � � �    X �      �    [ �  �������������?����������������� ��x�����������  xx������������0� �????��������	����������������8�8�8�p�������������������     � � ������          ������  ?00�z�f�    ???? � �������������    ������������ � ���'�8�g�/       ? ? � � � � ��� � � � �     � � � �       �����             � �����~�~        � � � ����6���6� 9 0   ��   �<�~�>�� ���  � �  ?    ��?��A�c�?`8�������������������������������������������                ��?��������    ??�������� ��6�>���������????��������q���� 7`a����������������~�����C�G��������������������W���� � � �����������������������������������������������ρ������������������������o������� � � � � � � � ��������� �`�`�� � � � � � � � �    ?.�.��         ?  6�1�g�'�?����  � �  ? ? � � ���0�� � � �    � � � � � � � � � �             ?  � � � � � �>          �����������������#i`���������������������                 ��������~��� ���������  �� ������������������������A�$�|'���������������������� �!�c ���    ����������������'�#�m���   ������������������?�h8�0�`�`   �����������������@�@|�\������������������1s{ x 0        � � � � � � � ��8�8�8� p p `    � � � � � � � ��@'� �v v r `    � � � � � � � �� @�G g � `      � � � � � � � ���?pq� � � � � ���>>  	y � � � � � ���   	����.;�l�~�w��H�<   �      � � ��;�3�wX��|�~p��   8 X     p �                               �<�����    ??����x�8�<�<�8�x������������������ � �           ����������������          ?                        � � � �                ���<�x������������������������<�|�������������������                 � � � � � � � �                 � � � � � � � � 		  � ���� � � � xp��������x� � � ���        ���� � � � ��� �        &2 p � � � � �          � � � � � � � �? ? ?     =  � � � � � � � � ?���>�>�  ????������(�������������������� � �Ќ � � � � ����������������                ����������������?�?�0�p�`�����??????���������������8�8������������������</?�!�7������������������<�|�x�����������������������;�l�~�w��H�<   �      � � �          � � � � � � � �        ?                 �`�0�0          ``0088 ��������������  ����������1�(� �$�,�>�B���????????��  8 >731         0� ~ < | � � � �00      w�|``000� �  ����������88  �F� �  � �??          ��������������pp!  � �N�.�<�L���İ��88    � � �      ?c��A� �     99qqAA��������   �������� ��� �`�`_���� � � � � � � � �-�!�p�0�O��3��  ? ?  ?  � � �  < ~ ~ �8�8�8�  88888888 s1�{�{����w�              ��`� � �` � σL                 ?   � ��?<<        �� ~ � � � � � � �8800      <<<<    � �gc1         88��/�g�s�/���     ``p      �p�p������t�p�     ���     � � � �� ��         � �  ? ��	��        ��0���o�?�Oy�{� � � � � � �    ��0 � � �@���?         � x <  �                       � � ���0�3�         ? ?���&�<�$��8�    � � � � ���?pq� � � � � ���>>  	y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	            ���� �`�p`� � �  �   @ ` � � � 				             ����� @`�� �� ` ` ` @ �     �3 � �� �  � ��                 �3                       �  � �� �  � ��3                       �3                                       �@                                                       @�                �3 � �� �  � ��                 �3                       �  � �� �  � ��3                       �3                                � � � � � � � �                 � � � � � � �                                           � � � � � � � �                 � � � � � � � �                 � � � � � � � �                            0@ �                           ?  �&��>���    ? 9 1 3    � � �~�������?    � � � � � � & @@ @  @ @                   ��~�                   ? A>9
-U"�@@                 �  � �� �  � ��                 �f                               (((8d8D8D8d        (   8                 � � � | 8                                                                                       �                               � � � � � � � �                 � � � � � � � �    @@ @  � � ��                            |�0�            8 \ ����?�1� u    ? 1    �G~�|ψ�� �s� � � � � �   �                          ������?�?�                ������������                � � � � � � � �                                          ��������?                                                     ? ?  �                  � � � � � � �  �@��Ѐ�@� 0 �    � � � � �                       ? ?                     � � � � � � �           @�                 0�H� � |        | | 8            � ��|��o>�<�x�    � � o � � �  � ����    � � � � � �    >>~|�                �������?�                ����������������                � � � |�~�~�?�?�                   ? ? ~~�                �?�������                    ?�       � ����x�p�B�<�    ??����������� � �0� � �1�;�������??��   � x�t�� �x�x���������������� | � � � p    ����������������          @ � � ����������������                ����������������                ����������������  � � � � �???88 � � � � ����������}}���������� ?	�      	  ��������\����   ���\ � � � � �3����?�������{x   ��   8����������<�����?����{�?���}��x��������  } �� ���������|�<p��?�����s8�?�?�?�<� � � �????????<<      ��������� ? ������    z�@� ������� �����������ᇇ�����:��?�~������������ � � �8�x�p� ������������������ �          ����������������                ����������������                ����������������� � � � � �00       � � � � �   ���憆      /�6�8�>�<� � � �/ 6088>><<      ������c��� ? � ��g    ?�>�����������������������\��<����������������?�<�?�?�?�~�p� ������������������x�������      ���������� 0 8>>44>8    <<<<>>>>       >~8�x���        88xx���8�?�?�<�0� � �??????<<00    �1�����0�Z����������휜>>~~�����8�0� ��p����������珏<< ?  � � � � �����������������    ?�            ��;�bظƀ��� �  ����ww�;��� �8�<�~�F�$�>�6����Ø�~ V => ��   � x�t�� �x�x���������������� | ���_??����������������       � ��������������?���8� ��=�?���>>   = ?   ������������?���������8�0���o7�w������������70wpsp`o�����i��^����o��i� ^ �  ?��|�x�}}}}���� � �����?����    ��������O?      �� �������� � �������������    0�4�`���`���<<<<xxyyyy``�<�|�z�w��������������������
??  � �        L���l��;�3�  o��m;;33    H�@�������� ��������������5�7��������������7�����##���8�x�p� ����������������������        �?�???����������?�?�??  ? ? ?       ��?�������� � � � ����     1�s�c������������������������������`������ � �cc������������^�>�<�����������������?�����.����������??<< � � � �!�8� ��    9999;;?? � �p�������� �    pp��������  | �"�&�<�<�????>><<<<�>�<� �0� �������<<  00ppxxxx    ��y             �q��������  ������ ��~�b�%>6  ~ j => 6 �1����������8�??���������ޞ�>>�8�0� ��m-��~�����������-! ~ <�����f�}�m������� ~ }m� � � � �`��>�����������������                ����������������� ��>�>�?��x> > ?   �>���������~p������ � � �p �8� � � � � � p ���������������� �6ɼC�?  3c  66��������������[������||yy{{??����������������� ������������  ��=               �x�`������� � �xxxxxx������      ;>  �        �������?� � �����������     gO?        �� ���� � � � 1���ܜ���    c�3�>�6��������k ���������������z�w����������������� � � �`�`�������������������     ;�������������������=z?�?��?  = ? ?        �>�~�������� � �� � � �� �           8 x p   ������������������ �a#� � � �����������������~��\��������������������� ���� ��^������ᇇ���� ��������<�8�0�  ���ܜ�������  � �8����� ��      88����  ��� � �3����?�������{x   ����@����������<�����?������� � � ��#�!!���� 0� ��N��x�x����11�������� � � � ��??      �6�0�����H�|�l�����0 � � x | l                     �`������� �  ~~��������� � �0� � �1�;�������??��� � � ��� �x�x����������������             �����������������    ? ? ? >  ����������������!{.    �����������������#�s � ���� � ���������������� �B��aGG� �KKHH������##  �� � � � � � �������          ?�>�����������������������\��<����������������?r�@� ������� �����������ᇇ�����:��?�~������������???~ |              �|�,�,�||  ||<<<<      9                        �`�`����� � � �pp��������      z�@� ������� �����������ᇇ�����:��?�~������������� �B�$���$�B�  �B�$���$�B� �� �B�$���$�B�  �B�$���$�B� � � � � � C C c g    ` 8 < <    >�~���           ` p �  � � � � � ��                    ? �~�����                 ���p�p���������                                                ����8@8�8�8�8 � � � ��@ � � �                                ���� ���           � �����?� ���      ) � � �B�$���$�B�  �B�$���$�B� � ��8����<� �                 ��8����<� �                 �|����0�~� �                � �B�$���$�B�  �B�$���$�B� �� �B�$���$�B�  �B�$���$�B� � w ?80``��              ��?��@� �`����`         ` � � �ߏ��y� �� `           ������� � � � �       0    ���������?          � � �    � � � �������                �8�8�0�0@0@8�8� � � � ��@�@ � �                                ����8�p�p'�7�w    � � �   0 � ��x�0� � �x���          0 � � �B�$���$�B�  �B�$���$�B� � ��8����<� �                 ��8����<� �                 �|��<���|� �                                               = =    �         < < '�O�_���� � �  @ @ @ @ � @ p ��� �@�0� �0 � ��             � ��4�8�0�P���               ��y�?��������        � � � ? � � � <���       � � �   �� � �         �                �������� � � � � � � � �   = =    �         < < � �B�$���$�B�  �B�$���$�B� �� �B�$���$�B�  �B�$���$�B� ��`�8�0�?� � � �         ? 0?     � �  � � � �   � � � �B�$���$�B�  �B�$���$�B� �� �B�$���$�B�  �B�$���$�B� �    7 # c a �           > � � � � � � � �> ~ ~ ~ ~ | | }  ��$�� �  �   ~ <@y s��� �  ����� �� �   � � �� ?A?�?��a��w � �     � � �     ��O�G��p�� �               ~g�'��? � ��              � � ������� � �                ����<�8�p�q� � � � � � ��  � � ���?�#����> ~       � � � �B�$���$�B�  �B�$���$�B� �� �B�$���$�B�  �B�$���$�B� � � ����� � �   � � � � �      � � � � ��� �   @  0 �� �B�$���$�B�  �B�$���$�B� �� �B�$���$�B�  �B�$���$�B� � � � � � � � � � > ? ?     > � � � � � � � �Z!&   x x�>���~�>��?�              �8�|�~��A������          � � �  � � � � C C c a      8 < <   |#�b���`�    `�� ` ��? ��?�?�?�� � �                � ��x��                �?�>�>���@� �          @  ����`�q���� �� � @          0�`�`�`� 1{ � � � � � ��� � ���?�"���^�         � P  �����;��}�        �      ��0����g��|�            � ` ����8@8�8�8�8 � � � ��@ � � � ??                 � � � � �ppp < <             ?  y � � � � � � � �  ���>A� � �        �       x��|�|�8� ~ � �           �    aaa1qx0�8�      3 = @�A��� � � ��@ @            ������� �            |�|��G�?���0 �              � � � � ��p�p�p < <    � � � �      ?  y �  � � � � � �  ?�?���~�<À�=          � �^���ϸG��x� �P � �        }��?�:�����     � � � @ |����������:` � �          �8�9�7�?@���� � � � � @     �?�����������             p�����<�=�       < = � � ���|���         | � �  ?      � � � � � � � �   ���|<     �p�0� �0�P�A�!�����= } } y y � q s �#�C<�<�,SL� `����������?@?�9�8�8 ��� ��@��� �     ��� � � �     � ������<�=�       < = � � ���|���         | � ��0�0�`�`�`�p�p�p � � � � � � � �                                ��`b�7��~�              ��F�~�~��À��        @ � � ` ��?��8@8�8�8�9 � � � ��@ � � ��� � �  <x�?�            ?���q�0�0�� ?   q p p p �����p �       � � � �         �      � � �    � � �      ���8�� s   � � �  ��$�D� ������g o ~ | y � � � ����G�����  ���� �8�8�<�<@>@;�;������@�@ � � ?      � �� � � � � � x   ?���|�8�0�� ?   | x p p ����< � �       � � �          �0�0�0�0�0�0�0�0 � � � � � � � �                                ~�~�<�  ?                     x���p� � �    �               �;�?�?�?C?�?� � � � �� �@ � �~����������� � �                              
  
       �   � @ � @ � U � U � U * U * U � U � U � U � U � U � U � U �   �   � @ � @ �                                                 ��������||||||||������������������������������������������������                                          @ � @ � P � P �  *  *  
  
 U � U � U � U � U � U � U � U � @ � @ � P � P �                                                 >>>>>>>>������������������������������������������������                � � � � � � � �                 

��������@���@�����������UjUjU���U���U���U���U���U���U���U�����������@���@���                 � � � � | | | |         � � � � � � � � � � � � � � � � � � � � � � � �                � � � � � � � �                 `��`��P��P��5?*?5?*?U���U���U���U���U���U���U���U���`��`��P��P��                 > > > >             � � � � � � � � � � � � � � � � � � � � � � � �                	                        � � � � | | | |         � � � � � � � � � � � � � � � � � � � � � � � �                 

 � � � ��@ ��@ �*�U�*�U�*Uj*Uj�UU��UU��UU��UU��UT��UT��UU��UU� � � � ��@ ��@ �                 @@�@� p p   8                                > > > >             � � � � � � � � � � � � � � � � � � � � � � � �                       �`@��`@��P@��P@�
5*
5*

�UU��UU��UU��UU��UU��UU��UU��UU��`@��`@��P@��P@�                <~>~??    6ai�?�?�?�    � � � � � `���������                `�0����������                h0X0T8D8$$<                                  ������������������������                *�U�*�U�*Uj*Ujfffv333;p�p�p�0�8�8�8��          �@� � � � � |                             <��@� � � � 0                      62;      � � � `�`�                ����������������????????                
5*
5*

(8��(8                   (8Tl8�Tl(8                                                                                                 ��`�p�0�0�8���                            ���?������������������_���J� � �����������?��������                                                    (8                                                            ??������      ����?�����8�0�0�p�`���                                }�x�=����?����������������������?�����������?������?  l|                     8(��8(                     l|                   �B�$���$�B� � � � � �������?�� ���/�� � ����������� ����������������?�?������������?�w� � @ `     0                              (8                      (8��(8   (8Tl8�Tl(8                    8(��8(    �B�$���$�B� �������?�?���������?������������������3�n����7�g���������?�?�?��� ������s�����0�                                   ? _ ow{}~   ��<��Á���    ��<��Á���  ~xppppppx~� � � � � � � � � � � � � � � � �    � �|�8�� ?�?�?������/���������������������������0�b����������� ?)>P���7�y���`�`��1>!>��`�0���p�p���� �B�$���$�B� �~xppppppx~� � � � � � � � � � � � � � � � ~xppppppx~� � � � � � � �   ������<�� �    ������<���  ��?�?�?�������>�|����`� ���� ��0�a�C���|��Gx����9�|��?�?����?�{����.�\ܤ�l|9>8???�p�x��&�\ܤ�L| �B�$���$�B� ��>YySs##&���������i��x�x� � � � � � � � � � � � � � | 2       3?1?47| � �        f f                   ? 1           � � � �     &>����"#DG�ψ�HO���
�
�3���	�� � � � � �     � � ?     1 � � � � � � � � � � � � � � � � ��9�x�1������,������@�� � � � � �           f f   pw������`�`��g�g`�`� � �                                                     	   ������hx11�������������	��Æ � � � � � � �     � �       � � � �      � � � f f    � � � �B�a�a�Q�Q� � � � � � �<�b� � � � � � �!�A� � � ������ � � � � � ���� � � � � � ���&� � � � ��@���(� � � � � � ���L� � � � � �p����� � � � � � �� � � � � � � ���@� � � � � � ���L� � � � � � �8�E� � � � � � ���� � � � � � � � � � � � � � � � �I�I�E�C� � � � �A�A�#�� � � � �I�I�[�6� � � � ����� � � � ���6��� � � � ����!������ �h������ �`��� �D�D�D�B� � � � �x����x� � � � ���	�� � � � �@�����`� � � � �D�D�D�B� � � � �������x� � � � �$�$�l��� � � � � � � � � � � � � � � � � � � � � � � � � � ��� � � ����9�f� � � � � ��B�b� � � � � � ��"� � � � � � ���L� � � � �� ��� � � � � � � ����� � � � � � ���d� � � � � � �p��� � � ����?�� � � � � � �<�b� � � � � � �\�2� � � � ����� � � ������� � � � � � ���$� � � � � � ���@�:�D�N�;� � � � �B�B�F�;� � � � �$�4��� � � � �~�@�b�<� � � � �D�D�D�B� � � � � � �2�� � � � �������z� � � � �E�A�A�@� � � � ��� ����� � � � ����� � � � �A�A�#�� � � � �"� � � � � � � ����� � � � ���$��� � � � �/�H�L�'� � � � ��� �@��� � � � � � � �A�C�&��� � � � � � �<�b� � � � � �8�D�`� � � �@� � �.�1� � � � � � �A�B� � � � � ����,� � � � � � ��� � � � � � � �8�� � � � � � ���L� � � ����r��� � � ������ � � � � � ��� � � � ������F� � � � � � ���$� � � � � � � � � � � � � � � � ����� � � � �A�A�#�� � � � �<��B�<� � � � �!�"�"�!� � � � �G�D�f�3� � � � ��� �(��� � � � �����@��� � � � �t�����v� � � � �D�D�D�B� � � � �������v� � � � ����� � � � �'�(�i��� � � � �D�����k� � � � �$�"�b������ �@�@����� � � � � � � � � � � � � � � � �!�s�U�I� � � � � � ��� � � � � � �\�2� � � � �@� ����� � � � � � ���@� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �A�A�A�!� � � � �:�D�N�;� � � � �"� � � � � � � �������c� � � � � � �`���� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````````+++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�++++�++++�+++�+�+++��++++�+++�+����++�++++�+++�+��++�������+�+���������+�������������������+�������������������������������������������D�D������DD�D�D����D�D��D�����D�D�����DD�D�A�AD�D���D�D��D�D�A�AD�D���D�D�����A�A�A�A���A�A������A���A�A�A�A���A�A������A����A��A���A�����+������A��A���A�����+���A�++++�+++�+�++�A��++++�+++�+�++�A���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�j�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�*�j�j�*�*�*�*�*�*�*�j�*�*�*�*�*�*�*�*�j�*�*�*�*�*�*�*�*�*�*�*�j�j�j�j�ꢪ*�*�*�j�j�*�*�*�*�*�*�j�j�j�*�*�*�*�*�*�*�*�*�*�j�j�*����*��*���*�*�j�j�*�*�*�*�*�j�j�j�j�*�*�*�*�*�*�*�*�*�j�j�j�*�*�j�*�*�*�*�j�*�����*�*�*�j�j�j�j�j�*�*�*�*�*�*�*�*�*�j���*�*�j쪢����*�j�*�j��j�*�*�����j�j�8�8�8�*�*���*�*�*�j�*������*�*�j�*�*�*�j�j�*�*�j���*�*�*�j��j�8�8쪈���*�j�*�j�j�*�j�j���8�*�j��誢j�*���*�*�j��j�*�*�*������8�*�*���j�*�*�j�j�*��j�j�8�8�8�*�*�j�*�*�ꈪ�*����8�*�*�*�j�j�8�*�*�*�j�j�*��j�8�*�j�8�8�8�8�*�j�j�*�*�j�*�*�j���8�8�*�*�j�8�8�8�*�*�j�8�*�*���8�8�8�8�8�8�8�8�8�8�8�8�*�*�*�j�j�8�8�8�8�8�8�8�8�8�8�8�8�*�*�j�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8sss s�8???�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8�8{{{�x�x�x�x&s$s"s@s ?"?$?&?�8�8�8�8�8�8�x�x�x�x�x+++�8�8�8&{${"{ {�x333�8Bs`s@?B?�8�8�8�8�8�8�8�8sss�x 3"+$+&+�8�8�8�8�xB{@{ 3"3$3&3�8�8s`3333�8�8�8�8�8�8&s$s"s s@3B3�x�x�8kkk�8�x`s@3B3�8�8�8�8s(3"3$3&3�������X�xBs@s`3�x�X�X�&k$k
;;;s`3��{{{({H3B3�����������X`sJ?L?� ;";,;&;D3F33�8&{${"{H{h3������������x{j?l?&$" @?B?`s(3d3f3&3�8�8�8B{hsJ?L?�����ssssj3???B@`3�sH3b3N3{{�8�8�8FsDsl?&$" �;;;&s$s"s(s(?"?$?&?�`sJ?L?s`3sn3${
???{fsds s��B@ ;";$;&;��BsHsH?B?��LsJsj?l?s3sJ?L?"?$?&?&{                                                                                      l � �z�������~�]  $H|�������\]�l � �z�������~�]  $H|�������\]�      � ��� � �         � @ �@�        | �`� �           px                        p h �@� R r       0p<@,                            ���t�p�x�|�y�9��p`xppx{|}y{99  � �`�0�� ����    @` 0����~ H * � ��@  #   �   ����X~ H * � ��@  #   �   ����X.U*U*U*..��        . _  ~��H�@�@Ҡ�`��*�8   \@��l � � l � �z�������~�]  $H|�������\]�      � ��� � �         � @ �@�? ? ? ?          ����&�a�>��.�?�o��� ����&�a�>��.�?�o��� � �@�@0�P�� � @�H�� �        @        a �@� �         `p  	-og���O  ???8 d �@� D H H 0    8p 8 0 0                                   8/1        8;        ��,��`�       $����        ~ H * � ��@  #   �   ����X~ H * � ��@  #   �   ����X�O00 | <        /      � � q q � � � � ,  � � � � �                 < ^0�x�x�0~ <                       �  ��             @@        8 L0�x�x�0� | 8                 



� �B�$���$�B�   BB$$$$BB  � �B�$���$�B�   BB$$$$BB  � �B�$���$�B�   BB$$$$BB  � �B�$���$�B�   BB$$$$BB    � � ����    ? ? ~ ~ | | � � � � �� � �    � � � � | | � � � � �� � �    � � � � | | � � � � � � ��    � � � � | |  ~�{                   "                      � �`�|b            |   p h0X0\8,$        0 8                        < �<<��                        c�cc��                       ((((((((                



� �B�$���$�B�   BB$$$$BB  � �B�$���$�B�   BB$$$$BB  � �B�$���$�B�   BB$$$$BB  � �B�$���$�B�   BB$$$$BB  ���P�P�?�?  8@8@@/@/? ?      � ������ � 8 8  � �� �      � ������ � 8 8  � �� �     ������� � 88��� �      	                                   �:� ����    8 zssc   � ����{�wP/��    � � x p ��   ??����    ?   � ����������������� � � � � � � � �                                                � � � �                            BB<<<<<<<<BB     B < < < < B        @@    ��        @     ���         �                             > >        6> >               ~ _  /?  _ ~           ~ ^ ~ o  _ ~    0 ,      | �8�z�F���0<   8zF8bb<  p �p�@� �    p @0 `     p �P�Pp    
    P P            P                            ����?? � �   ?   ���������������� � � � � � � � �                       ? �                 � � � � � � � �    $$$$         $   $    ��ff~~<<<<~~ff�� � f ~ < < ~ f �      @@           @                          88TT������<<((   8 T � � � < (  $$  ��  ��  $$ $   �   �    $    � �B� � � �       1 I q A       � � � � � �       �           			           � �  �`�p�p     �   @ ` � � � ~ � � �� � � ~    f , f f    < < � � � � < <     ~ ~                      � � @�� � � � @   �   � � � � �         ? }� �\            ?          � 0              @��                                  ` � ��`            ��`` � ����P�?   ? ~ | 8@@/?   � � � � ����   � � | 8  ��    =ys�� �       A I Y � ��� � � � � �   ����$ � � � �                  ??������������  ? � � � � � �	             0�p�p�`�`@��� � @       �                      � � � � � � � �   � � � � � 0                    @ @ @ @ @ ����� � � � � �       �N � �7\?? ?    70?#     � � = ?���� 0�8� � ���   ��l�o67       llo'6         <�h����       ��hH��        � �B�$���$�B�   BB$$$$BB    ��||88llDD      � | 8 l D  � � � ^ S ;  Y Y I ) ,      � � = . j ����� � � � � �       ????������ ? ?    � � ����������������� � � � � � � � �< f � � � � f < < f � � � � f <   $ $ B B � �   $ $ B B � � � �PQ

         �P
          � @� @ ��DH         � @� @ 81          � � � �����  � � ` ``� �    <=              � � � H����    � � p  00�0          x              8         � x�4��          ` 8    8|6�>�>��   6>>wl` � < :$rL��✁�   @ �$�L�� �@�  !@?@?�I�I�I�            � � ����ܸ�|�  � | p ��������  / � �          /   @ � � � � � � �     � � � � �  � � � � � � � � � � � � � � � �     � � � � � �       �    2                                   $(	
	
         ! 8<          \����0�� � � 0�`�� � �   sC<A>8   3       ������0�� �� � 0�� � �   |���~�b@ > < y s  ?    ������|�� � �� �� �   I9�g�ow?  9go       ��b���� |�� � � b�� �   �     �~?|7!> 8? ??77      |�� � � < ~  � ��x X � � � �   |� o �/  0 0          ���� 80��� @ �8 � � �                          p�p �          P                ~ �~�~�             ~  � � � | ?      ` p 8       /+/'          � 0�� � Ԁt ��   @ � � x � � �   @&@ �H�@                � 0�0                      @&�F�P                    � �                                    �  �                   9yk�0�0�     0 " F O  � � ������  � � � � � � �                                        � � �             � �  @#@'@'�O�O�O�G               � � � � � �                     $f$�Z�[f$$ < ~ ��$�$�~ <      <<          < <      ?:/.              ��(�H���0��� � � � � � �     �@�@@ @                   "$00��                �@�@@                       "$��                                        $(HP  ��        @        � �  @     o O 0 ?       ��<8����� p 0 � � �       >>               � � � � � 0 �08 � @ x � ` �            $                     < ^ f f z<                      <f$f$<      < ff<                                 �������G  < | ~ ~ ~ | 8 � �������    < < <  3gN1�"�@�@      � 8��0�����       ����������� � � � � � � �          � � � � � � � �   � � � � � � �     ` �`�p�pL0J4                 $$&I6I6�l�                         ?                   � � � � � �                  <B=�x�p�c`'p        @ � ��0���     � �p0p  @8`0p�;�           � ��,��      � �00�p �p�xa@?I68                 ` �`�`H0H0�x�\a                ���x�p�p�p�?       O@08   ���~~y~�� <   ���x�   �@�p�0O0o0           � �3��<0��� ������ 0��   !!    ��!!    ��� � � � � � � �     @ ` � � � � R,B<F8I6�~�l�``                 		`�|�nn                 ?    � � � �                 � � � � � � � �                 �~�|�~�L48  @@` 4   ���np�� p ��  ��| � p  �~�~�N>6  @` >    |��s|Gx>�� � �� ��~�~ � �        � ���p�                  ���p�x�l�ny                                                                              ~~����~~xx��cc  ~ � � ~ x � c77������   7  � � � ���������������� � � � � � � � �00yy{{kk    0 y { k �����������ޞ� � � �  � � � �      00            0             ��          �   qr���p�``    0 d h        0@0�c�g�           @� x�$���      � �8� 9 %"0            � �\���pp ����    � � p� @ @ ? oP?W8T8W8_?`         � ����8T8�8���  � �    � �   <<~~~~<<  ��     < ~ ~ <   �    <<  @@      <    @     ll������8888   l � � � 8 8 ������?????? � � �  ? ? ? ���������������� � � � � � � � �����qq##99 � � q #  9  TT����^^LL����   T � � ^ L � �      !!           !        ��  ��      �     �    < B<�v�b�B�fB<<                 �~` `?r>_?# `    2 ?   ~~��4848�� ��� ��8�8 �               ��������� H  � @ @ @ @   ����  ?            � @�x�h�x�h�H��   � � � � � �     ?~   >� � ��������w��t  � ���𸻹�pv�        � � � �@               @�����t�p�x�|�y�9��� xppx{|}y{99  � �`�0�� ����    @` 0����      ?         6� � �� ����   � 0�0�����         � � � @                �                       u������� � �hP"��aziL N��  � ���������    @� ���� �������������   ������������� ���`�������   �F`������     ?~         >� � ����������   �����������       � ��  � �          �@�   `� � � �x0  ~G8~ 8     �8�=�}<��s��t�z�~�<�<<  x@| � � � � @ �      @`      �      8??;c>G> 8;  $8   ��(� �x�x^��� $��  ```��  ����3 .nnO.w;    � � ����>�� �� � � 8     � � � � �   @��                                        �?�� 3c?G?    $8   �p��� � ��|�|� �|����pp  ` p   �<�0?? c<G> |}>>?   $8   ��� �x�x^��� ��  ```��  ����y0 {{C;}8     ������������:�0������������ >0� � � �   � @ � `0@   @ �   �     ?       ` � �����������   @���𰴰���      ?     (� � �� �0� � �   ` `� ��0�0� �    �� �      ��� ~�~��"�B� �0�0  �(�(&*BB82�2��8�=�}<�Y�S����~�<�<   `    ����� �0     �g205x  � �������>��    n���~��>��  � � �1�!�   3 	05y%yM1� ��8�x��������  8�8�x��������                         u�����0�0� � �@P"�� =2|6x>@< A@  � ���������    @� ���������t�p�~���?��� xqp~~??x � � � � ������   8$�L�| ������    < 5 ? ?#?      ����~�?�6��8~�~���00����x& PPPn 0     �� ��9�*�,������ �     �����x�0? G> ����?      � � � �`�x^��� 8�   ```��  �8�=�=<�9�s��4�z�~�<�<  8 | �!�  ;c?G> %yM19 $8   ����� � ��|�|� �������� ` p   �� ? 3c?G> ;??   $8   ����� ���|�|� ������@@ ` p   �8�=�}<�M��� �~�<�<00a  �`�?`??    �p��� � ��|�|�8�|����pp      ( ??? 	??      ����� ���<�|�x�8������� 0 p `0                     0   ���    0 ????�����������  0   ����������������      ������ @p0      ����������zd{dwhsLgXC|��{~������=��?�C;��������������{{�|�x��L���w{������������������:4���¦�{=�����������������  @�??���   " 0a����������������""���ޜ�99##GG""���ޜ�99##GG����pw &���ܱ�xx����ww&&���ܱ�xx��������??~�nn��������??��nn��������������??��������������??? 3GxmS@?��????�����`�0��|���<���������������� 	p � � ? <@p�`����������������� � � � � ? s�<����������������P0`  P  ����������������~��	����;;�~~������������3{������ߜ�33{{�������ߜ�����0���8>p��������>>���c	� �x0^`��������~~??~~��FaLc��������������������$� ����V^}}pprr��������^^}}pprr@@�Ο�SS&&  @@�Ο�SS&&  ````      ````      ppccGGFF������ppccGGFF������??��33<<88??��33<<88����;���������@@��������������@@r�������������������������������                    0   ���    0 ????�����������  0   ����������������      ������ @p0      ����������zd{dwhsLgXC|��{~������=��?�C;��������������{{�|�x��L���w{������������������:4���¦�{=�����������������  @�??���   " 0a����������������""���ޜ�99##GG""���ޜ�99##GG����pw &���ܱ�xx����ww&&���ܱ�xx��������??~�nn��������??��nn��������������??��������������??? 3GxmS@?��????�����`�0��|���<���������������� 	p � � ? <@p�`����������������� � � � � ? s�<����������������P0`  P  ����������������~��	����;;�~~������������3{������ߜ�33{{�������ߜ�����0���8>p��������>>���c	� �x0^`��������~~??~~��FaLc��������������������$� ����V^}}pprr��������^^}}pprr@@�Ο�SS&&  @@�Ο�SS&&  ````      ````      ppccGGFF������ppccGGFF������??��33<<88??��33<<88����;���������@@��������������@@r�������������������������������                    0   ���    0 ????�����������  0   ����������������      ������ @p0      ����������zd{dwhsLgXC|��{~������=��?�C;��������������{{�|�x��L���w{������������������:4���¦�{=�����������������  @�??���   " 0a����������������""���ޜ�99##GG""���ޜ�99##GG����pw &���ܱ�xx����ww&&���ܱ�xx��������??~�nn��������??��nn��������������??��������������??? 3GxmS@?��????�����`�0��|���<���������������� 	p � � ? <@p�`����������������� � � � � ? s�<����������������P0`  P  ����������������~��	����;;�~~������������3{������ߜ�33{{�������ߜ�����0���8>p��������>>���c	� �x0^`��������~~??~~��FaLc��������������������$� ����V^}}pprr��������^^}}pprr@@�Ο�SS&&  @@�Ο�SS&&  ````      ````      ppccGGFF������ppccGGFF������??��33<<88??��33<<88����;���������@@��������������@@r�������������������������������                    0   ���    0 ????�����������  0   ����������������      ������ @p0      ����������zd{dwhsLgXC|��{~������=��?�C;��������������{{�|�x��L���w{������������������:4���¦�{=�����������������  @�??���   " 0a����������������""���ޜ�99##GG""���ޜ�99##GG����pw &���ܱ�xx����ww&&���ܱ�xx��������??~�nn��������??��nn��������������??��������������??? 3GxmS@?��????�����`�0��|���<���������������� 	p � � ? <@p�`����������������� � � � � ? s�<����������������P0`  P  ����������������~��	����;;�~~������������3{������ߜ�33{{�������ߜ�����0���8>p��������>>���c	� �x0^`��������~~??~~��FaLc��������������������$� ����V^}}pprr��������^^}}pprr@@�Ο�SS&&  @@�Ο�SS&&  ````      ````      ppccGGFF������ppccGGFF������??��33<<88??��33<<88����;���������@@��������������@@r�������������������������������                      � �(   � � � � � � �      7        ?         @�P��$�   � � � � � � �                 $ $ <       ~~<<<<ff   $ � � B B � �              <          ����������    � @ @ <     ??    � � @     ��������������� @ `   ?                                     B < < < < B                  � � � � � � � �  � � � � � � � �� � � � � � � �  � � � � � � � �� � � � ? � � �  � � � � � � � �� � � � � �  /  � � � � � � � � `       � �      �$��� �  �`   � � � � � � � �<$          ?      � �  �      � � � � � � �       8             8         �         �                    ������pp         � h      88         ! F X ` ��������xx      � b        $   $                     � f ~ < < ~ f �                � � � � � � � �  � � � � � � � �?    � � � �  � � � � � � � �� � � � � � � �  � � � � � � � � O  � � � � �  � � � � � � � �� � � � � � � �  � � � � � � � �� � � � � � � �  � � � � � � � �� � � � ? � � �  � � � � � � � �� � � � � �  /  � � � � � � � �� � � � � � � �  � � � � � � � �� � ?  �  ?   � � � � � � � �� � � � � � � �  � � � � � � � �� � � � � � � �  � � � � � � � �                     D (  ( D                       D (  ( D                       D (  ( D                       D (  ( D  � � � � � � � �  � � � � � � � �� � ?  �  ?   � � � � � � � �� � � � � � � �  � � � � � � � �� � � � � � � �  � � � � � � � �� � � � � � � �  � � � � � � � �?    � � � �  � � � � � � � �� � � � � � � �  � � � � � � � � O  � � � � �  � � � � � � � �� � � � � � � �  � � � � � � � � � � � � � � �  � � � � � � � �� � � � � �  �  � � � � � � � �� �  � � � � �  � � � � � � � �                     D (  ( D                       D (  ( D                       D (  ( D                       D (  ( D  � � � � � � � �  � � � � � � � � � � � � � � �  � � � � � � � �� � � � � �  �  � � � � � � � �� �  � � � � �  � � � � � � � �� � � � � ���� o`������������� ����� � �  ����{x�8�8wp��� ����� � � ����;8�8�8wp��� � ������� �0�0wpwpo`����� �������� � }|����? ����� � � � � � � ? � � �   ������  � ��8}\}}{x�8�  ��� � �����P� � �	���� � �  h��82� �� �������� ����������  � �����?�8�0� �� � g ����wp� � � ��8�<��� ��wpwpwp������ �?�?������ �������������� ��� � ���� wpwpwp������? � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �| ~Z Z Z Z Z Z Z Z  � � � � � � � �� � � ������ o`������ ����� �����3� � � � �;8��������� ������� ����=<�8wp����� ����8�8�<� ������wpwp����� ������� ����=<����8 � � � � � � � �� � � � � � � �  ������  � � �   ������    �     ������  < � � � � � � � � � � ���8�8�<��� {x�8�8wp������? �������� ������������  ���8�0�9��� �������������� �������� ����������  � ���8�8�<��� �8�8wpwp������?  � � � � � � � �  ������ ���  ����   ��U �    ����   ��U �    ����? ��`A�#�"Pp"Pp"Pp"Pp� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��	 ? ������������������ � � ����G`��'�0��  � � � � � � � �� � � � � � � � �
��
��
��
�� � � ������ � ? ���p����������� � � �������� � �  � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � �� �~�`�|�`�`�~� � �<�f�f�>��<� � � � � �<� � � � �<�f�f�~�f�f�                                                                                                                                                                              #                          0 �0�                                        � � � Հ׀�����@ 0@8@8 ( (   �@�@������������ 8   > 
       ` � � ����׀         ` p p (_ > >.&�@C�� >                     �p�                                                           0 �0                                                                                                                                                                                                   �? � � � � g             � � �� � � � � �              @ � �o�m�#�#@    0         �����@�������p� | 0        � ��������v���              �ց��ԃԃ����� � ( x ( ( 0     ? � ����@?@?@?           � �� ������ � �           #�?@�`� � ��g�             |�� � � ���`             @ �  ` �`��d�| �           �                                                                                                                                                                   � h             o               	 �   � � �       L0�|� � � � � �          0 �     �p� � ~ <�{�1� p     � �    � B�<��( ��<~ <    � �   �p� � � ���� p         � � � � � � � �                 � � � � � � � �                C Q ) &�"���� � � � A A a    � � � { 3   �        � � � � 7 � � � � � �               p � �                                                                                                                                                                                                                                 �          � �               , �        � � � �        (�    �        � � � � � � � �                 � � � � � � � �                 � � � � � � � �                ��������   0 0 0    4             �q� � � ��� � p            �����������������������������������������������������������������������������������������������������������������������������������֪�����V�VҖӖ���֨��ֺ�������ٖؖ���V�V�V�V���ֺ�����ᖹV�VÖ���ָ��֪�������Ȗɖ���V�V�V�V�����������������ٖؖ�V������V�V���֨��V�V����㖸������������Ȗɖ�㖸����㖷V�V���ָ��V����V�V���������V�V�V�V������ҖӖ�������V�V���������V�V�V�V���������V�V�V�V������Ö�������V�V����������V�V�������ְ������������������������������������֠�����������������������������������������������������������������������������������cd��������������������cd�����pqrst�����������������pqrst����fghijk��dUcU����������cdfghijk���uvwxyz{��tMsMrMqMpM����pqrstvwxyz{���lmnopFG��kMjMiMhMgMfMuM�fghijkmnopFG���|}~DEVW !{MzMyMxMwMvMlMuvwxyz{}~EMDMVW !"#$%TUP01GMFMAoMnMmM|MlmnopFG$%UMTMPP012345PPRS@AWMVMEMDM~M}MuM|}~EMDMVW4RSPPP@ABCRSPPPPRSMPMUMTM%M$M#M#~CUMTMSMRM5M4M - -b111 - - -L1M1 - - - - - - - - - - - - - - - - - - - - - - - -111111\1]1 - - - - - - - - - -MqLq
111 - - -L1M1 - -(1)1*1+1,1-1.1/1N1O1 - -MqLq11qqq
q]q\q111111\1]1 - -8191:1;1<1=1>1?1^1_1 - -]q\q11qqqqOqNq*1+1,1-1.1/1N1O1 - -H1I1J1;1[1[1[1;q&1'11 -OqNqN1O1-q,q+q*q_q^q:1;1<1=1>1?1^1_1 - -X1Y1Z1[1[1[1[1[1617111_q^q^1_1=q<q;q:q*1+1;1<1[1[1[1;q&1'11 -e1K1[1[1[1[1[1[1[1;q&1'1N1O1Y1Z1[1[1[1;1<q;1K1[1[1[1[1[1617111;1[1[1[1[1[1[1[1[1[16171^1_1K1[1[1[1[1[1[161[1[1[1[1[1[1[1;q&1'1��      � � ��                     88|8|0                ���{���o                �`�������������                ��	  &_ |~       0(  �+����� ��� �   @� �  ��� ����[� ? �  �    � ��m � �� �D�� � � � � � � � ������G �`� � �������    � �� � � � � �          ���� ,�? � � � � � � �         �? � � � � � � �              ���������000                � � � � � � � � ��       � � � � � � � � ���? ? ? ? ? ? ` ` @ � � � � ��V�V� p p �p�p��                �t���h|>>O>�                �V�Vs????�;                ����������������                ���xt����00 <<    0<������p�?�?     x00  ��� � �h�Z�9~�    hhXX8888@�G��@�@����~�|�� �   �����/`�p�p����0 0 ������ � � � � � � � �          �� � � � � � �                 � � � � � � � �         ? �������l �                 � � � � � � � � �� � ��� � � � �  ?    ������ � � � � �  c  ��� P Q                    >>���������                ����ߎ����;                ������� � ��Á                uM�����y�w��� <? ?   <�? �@�� ��p�8�0  ��@� �@� x 809lMu��w�o�W�;((hhpp``PP88����������������      |Ml�`�`�`�`�`�`����                     � � � � � � � � uM|          � � � � � � � �   �               � � � � � � � #M#� � � � � � � �                 � � � � � � � � � � � � � � � � ��               � � � � � � �  - -                     ����?�?����~ T               - -�����_��_                � � �����@��@�                 (1)1txtyw{< ??   �00�O���@���� 0�� ��� �   8191;�;�?����00 � � � � � ���������������@         A@H1I1�>� � ���  ? � �   � �o �	� ���@�� � � � � � � � X1Y1!� �� ��@�� � � � � � � �     � `�0�8�x�� � � ? � � � � � e1K1� � � � � � � �     0` �@��� � � � �  ? ? ;1[1 0          x � � � � � � �   � @   0 �  � � � � � �                                                � � � � � � � �           � � � � � � � �      A � �      � � � � � � C       � @      � � � | � � � �  c !   @      � � 1 # � G  |� � �            � � � � � �  <                � � � �  ? � � � �������������    ������������               �                        ?              � ��3�������      ??������   � � ���������        ��������                                                                                                              � � � � � � � �                  8 p �             p g � p  �      � p        8      z � �  8                                               � �   x a �       0 x � � �  � �  0 x � � �    X �      �    [ �  �������������?����������������� ��x�����������  xx������������0� �????��������	����������������8�8�8�p�������������������     � � ������          ������  ?00�z�f�    ???? � �������������    ������������ � ���'�8�g�/       ? ? � � � � ��� � � � �     � � � �       �����             � �����~�~        � � � ����6���6� 9 0   ��   �<�~�>�� ���  � �  ?    ��?��A�c�?`8�������������������������������������������                ��?��������    ??�������� ��6�>���������????��������q���� 7`a����������������~�����C�G��������������������W���� � � �����������������������������������������������ρ������������������������o������� � � � � � � � ��������� �`�`�� � � � � � � � �    ?.�.��         ?  6�1�g�'�?����  � �  ? ? � � ���0�� � � �    � � � � � � � � � �             ?  � � � � � �>          �����������������#i`���������������������                 ��������~��� ���������  �� ������������������������A�$�|'���������������������� �!�c ���    ����������������'�#�m���   ������������������?�h8�0�`�`   �����������������@�@|�\������������������1s{ x 0        � � � � � � � ��8�8�8� p p `    � � � � � � � ��@'� �v v r `    � � � � � � � �� @�G g � `      � � � � � � � ���?pq� � � � � ���>>  	y � � � � � ���   	����.;�l�~�w��H�<   �      � � ��;�3�wX��|�~p��   8 X     p �                               �<�����    ??����x�8�<�<�8�x������������������ � �           ����������������          ?                        � � � �                ���<�x������������������������<�|�������������������                 � � � � � � � �                 � � � � � � � � 		  � ���� � � � xp��������x� � � ���        ���� � � � ��� �        &2 p � � � � �          � � � � � � � �? ? ?     =  � � � � � � � � ?���>�>�  ????������(�������������������� � �Ќ � � � � ����������������                ����������������?�?�0�p�`�����??????���������������8�8������������������</?�!�7������������������<�|�x�����������������������;�l�~�w��H�<   �      � � �          � � � � � � � �        ?                 �`�0�0          ``0088 ��������������  ����������1�(� �$�,�>�B���????????��  8 >731         0� ~ < | � � � �00      w�|``000� �  ����������88  �F� �  � �??          ��������������pp!  � �N�.�<�L���İ��88    � � �      ?c��A� �     99qqAA��������   �������� ��� �`�`_���� � � � � � � � �-�!�p�0�O��3��  ? ?  ?  � � �  < ~ ~ �8�8�8�  88888888 s1�{�{����w�              ��`� � �` � σL                 ?   � ��?<<        �� ~ � � � � � � �8800      <<<<    � �gc1         88��/�g�s�/���     ``p      �p�p������t�p�     ���     � � � �� ��         � �  ? ��	��        ��0���o�?�Oy�{� � � � � � �    ��0 � � �@���?         � x <  �                       � � ���0�3�         ? ?���&�<�$��8�    � � � � ���?pq� � � � � ���>>  	y     ��(�           ? >  �������?�c�   �  �    � ��^�������� �    � � � � � �        � ����� �          �      ?s>�0� �h�X��     ? < 8 x x ���t����3 3   � � � <    �<�L���|�X�I�   ?  | | ?   �|��!�y�{ ��-�   � > ~ | � � �       0``                  ��p������         @ � � � � ��>�?���|�0       8 | x | 0       � ��<��                �`�`�a�g�g�g�   0 w g N  7 w � � � �������     � � � � � � �����{�����    � � r � � �f���=���� ��� � � � � �    �&�#|7xy{  => > ?        f�@� ��> ��,��0` �     | |��`� � � � � `� � x 0         d�|�<�,���.� � | | < > > > >  �`�`� �lx  x x | ?      s(�h���0�  8 �  < | � � � �  ��y� � � � � � O   q q c ,  ��3 7� � � � � � � �    ?X?��O��?`?�?�  8 0        � � � � � � ��              � � � � �����            ���?�����������  < | � � � � � � � �W�w�0� �  w w w w w s 0   � � ���    � � � � � � � �    
�����1 � � � � � � � �   \��?����|�?��� � �          ��?�?�?�?��  8 | ~ ~ ~ | 8  ��������      > > > ���?_???��� � � � � � �  ���������������� � � � � � � � �0� ��� �0�0�  ? ? ? ? ? ? ? ��3������  � � � � � � �0�?�����?�0� ? ? ? ? ? ? ? ?�0� � � � �0�� � � � � � � � �?�o ?                  ����<�8� �  ?  � � ? ?      ����<� � � � � � � � � � � �    �� � � � � � �   � � � � �       ? ? ������           0 0 � �� �� � � �      � �         � �8�p�� ` �        � �         � � ���      � �    �����?� �       @p8  ������ � �>   ���~ �  @� �0��� � � �? ?         �8��� > � � �� � � � �         8xw���        7 /  �����8�h8     > � �� �A>�`�@� ��p��  �  `@  @� �����g� ?  ` 0  x ���0�0�0�3�3�3�0�0� ? ? ? ? ? ? ? ?��3 � � � � ��3 � � � � � � � � � �`���������    � � � � � �   ?����������     c � � � � /�/�/�/�/���� 0 0 0 0 0 0 0 0� � � � � @ �                     ?78	17?              � ����8� �    � �  �          <?? ?               �?������      ?  � �  � � � � � � � �    � � � � � �   ? � �0�p���@�      � � � � �~�4� �a�c���' G  8 x|0 �<�x��������� �  < x���� ��?���������� � � � � � � � s,�<���������� < < � � ��  � � � � � �0�8� ? ? ? ? ? ? ?  � �����=��� � � � � � � � ?���� � � � �� � � � � � � � 
�������� 0 0 0 0 0 0 0 00`�             1 c �                 �0t����        ���?@?` 0<� � � � � � � � ??    �        p�p�l�h�x�x�@�@�L L |   < | |  � � � � � � � �� � � � � � � � 0�0�0������ ? ? ? ? ? ? ? ?>�>�<�x�p�4�$��    pp    � � ? ~ � ��������?o 0<� � � � � � � � �� ;;< x � � � �����/��� ? ? ?          �� ?�� � � �� � � �         �������� � � � � � � � � � � � ��� ? ?     0 8          <?y � �         ?     �  ?  ��� � �         � �    ������ � �    | � �    ��� � � x  ? ? ?         [�� �5�5� ��    [       [ ���� ����� ��   � �         �     <?? ?                �:�d�����      = { � � � �� � �   1 !          @��w �����/� �    , H �  ��� � � � � �`  �           `�x�v���h�4��� � � � � x <  �� ������    ? ? ? ? ����o���9g��w� � � � � � � � ���� �1�b��/���� � � � � � � � �    @��� � � � � � � � ����?��<�x�x� � ?   � � � �������~����� � � � � � � �                                                                 ��� �5�5� �� [ [ [       [��� ����� �� � � �         �
64y,s8g      < 8 p�`�a��3�0ϥ�L�� � � � 9 q � �             o _ � � �@�@�@�� �       @ @ @ @�@�@�@�@�@�@�@�@ @ @ @ @ @ @ @  � � � � � � � �                ��������? ?       ��������=�x�� � � � � � � � �����-��>������ � � � � � � �    �  � � � � � � � � � ��|�����9�@�� � � � �   8       ���� �         � �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   ���9��  ���=��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ^�6o^�of�of� oV�oV�oU�oomgm"o&m�+m �+m"g mu.m�z j��j��j��j��j��
j�b*�b*��d*�mi�eim&i��+i �+ie i�s.icc[cc&cy+cy+c[ ci.c$`a$Xa,`&a%v+a*v+a,X a#f.aH`eHXeP`&eIv+eNv+ePX eGf.edfgd^glf&ge|+gj|+gl^ gcl.g��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��         ��b�� ( 
               �_�g�1�-�6�W��%2[�  �%O�HA�!v!�!�-�6�W�1W6=S�w�!���#9g��yu�{����(�)�)d*�#�H1'e0S�[�g�g�R�c�k�s�{����#9g�Y9YB�J9K;�Q�Z�s�Q)�5_[�#��9�#�#�#�G��{���S�c�s��-9g�S9WB�J7K�1;�Q�������#9g�T]Xfg8g�1_�Q��0S�_�o�{�:     �� Fp ?'W�k�_Q  �AU=�$�eF �U�~?W�k��G  � e ��F �?W�k�k  �E� hb�F q�_?W�k�9~  
E$ qe�8F �}_a?W�k��  � �� F�?_'W�k��  nD%��iNF_!Ng?'W�k��1  B$�$ �@�8F k]_Q?W�k� �        �AA� � � � �   �                � p h      � � @  9K9�J  K  �� �A      N ���    �                        � �                           �   �   i A  l       ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    Q)�    Q)�    Q)�    Q)�    Q)�    ��    Q)�    Q)�    �5�    Q)�    Q)�    Q)�    �5�    _[�    Q)�    Q)�    Q)�    _[�    �5�    _[�    �5�    Q)�    Q)�    Q)�    _[�    _[�    ��    ��      �      �    Q)�    Q)�    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    Q)�    Q)�    Q)�    Q)�    Q)�    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    Q)�    �5�    ��    ��    ��    ��    Q)�    ��    �5�    �5�    �5�    �5�    Q)�    _[�    _[�    _[�    _[�    _[�    _[�    _[�    _[�    _[�    _[�    ��    ��    Q)�    ��    ��    ��    ��    �5�    Q)�    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��    ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      � �       ��     ��      � �     � � �   � �        � � �   � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        ^ � 6  ^ �   f �   f �    V �   V �   U �   p    h   " p &   � +    � +  " h    v . � {    � �   � �   � �    � �    � � 
  � � b   � � b    � � d   �n   �f    n &  �� +    � +   f   �t .  d    \    d &   z +   z +   \    j . $ a    $ Y    , a &   % w +   * w +   , Y    # g .  H a   H Y   P a &  I w +  N w +  P Y   G g . d g   d _   l g &  e } +  j } +  l _   c m . � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �        � �            ��������������������������������V   � ��^   � ��V 	  � ��^ 	  � ��V   � ��^   � ��W   � ��g   � ��_   � ��g   � ��_   � ��g   � ��_   � ��g   � ��_   � ��g   � ��_   � ��+   � ��#   � ��   � ��+   � ��   � ���   � ��*   � ��"   � ��h   � ��%   � ��b   � ��r   � ��b   � ��c   � ��c   � ��l   � ��t   � ����������������������������������������������၁���၁���������������������������������������������������������񱱱����������������������������������������������������������������ѱ����������������������������������������������������������������������������            e�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ���~�  ` *v��    `  !��  (  +$���
  (  +
���<   �  J���w#   < �PPw ��     , �����  � �R�\��4�����^  �~�� �ܢ�� ~ ���zު���^���x������6�O�  �    XF0X���
�	8�P��;L���   �.V�$&F��B�	��!c���  4	N�Fn�f���N�:N�9��� <  �x������ �.�)" ~P<��wo w  �   � �  �  � � ( ��@  �     �����  �z t�"�0�J��L)���  8����w��l\ ���&A�l���)�   @M�  �    �< ʢ��, C��C����H<� ��-                                                                                                                                ��G��������    1   �6    ��� �    � �6�  ���ݶ�             @�                        �6        ?g��:��<� �� $=�� �
����w>���?��t�Q��=�xܶܵ?����#?�+�
�>�e�#��=�=�J=�M$p���=�#>T�?iл:��<� =����ܲRf�b!>X<����=2">T�?b����
`��=8�ZT�jjdd
`�YSiicc
`=�V>f`�`=�=1�!>T>�<�������v�6�7�,=@�=I>`A>t�%P&P'P�c����=�� �x�rh>o�X=�x	'>��'%���`=�Z=@��Z=@PP>�=�M=�I�"Z�0�u=�� ePW�,�=>�1"R`>����?=�>!��
ӥ�ue	)>�>�>�=� >�=�>�>��W�� �==�uem!c>�.�M=�޵4��=ʶ4��=�,�!P)P*P��<,=��>`c=��=����@�P>��@���� �                         � d                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 